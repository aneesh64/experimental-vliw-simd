// Generator : SpinalHDL v1.10.2a    git head : a348a60b7e8b6a455c72e1536ec3d74a2ea16935
// Component : VliwSimdSoc_1c

`timescale 1ns/1ps

module VliwSimdSoc_1c (
  input  wire          io_csrAxi_aw_valid,
  output wire          io_csrAxi_aw_ready,
  input  wire [31:0]   io_csrAxi_aw_payload_addr,
  input  wire [2:0]    io_csrAxi_aw_payload_prot,
  input  wire          io_csrAxi_w_valid,
  output wire          io_csrAxi_w_ready,
  input  wire [31:0]   io_csrAxi_w_payload_data,
  input  wire [3:0]    io_csrAxi_w_payload_strb,
  output wire          io_csrAxi_b_valid,
  input  wire          io_csrAxi_b_ready,
  output wire [1:0]    io_csrAxi_b_payload_resp,
  input  wire          io_csrAxi_ar_valid,
  output wire          io_csrAxi_ar_ready,
  input  wire [31:0]   io_csrAxi_ar_payload_addr,
  input  wire [2:0]    io_csrAxi_ar_payload_prot,
  output wire          io_csrAxi_r_valid,
  input  wire          io_csrAxi_r_ready,
  output wire [31:0]   io_csrAxi_r_payload_data,
  output wire [1:0]    io_csrAxi_r_payload_resp,
  input  wire          io_imemAxi_aw_valid,
  output wire          io_imemAxi_aw_ready,
  input  wire [31:0]   io_imemAxi_aw_payload_addr,
  input  wire [2:0]    io_imemAxi_aw_payload_prot,
  input  wire          io_imemAxi_w_valid,
  output wire          io_imemAxi_w_ready,
  input  wire [31:0]   io_imemAxi_w_payload_data,
  input  wire [3:0]    io_imemAxi_w_payload_strb,
  output wire          io_imemAxi_b_valid,
  input  wire          io_imemAxi_b_ready,
  output wire [1:0]    io_imemAxi_b_payload_resp,
  input  wire          io_imemAxi_ar_valid,
  output wire          io_imemAxi_ar_ready,
  input  wire [31:0]   io_imemAxi_ar_payload_addr,
  input  wire [2:0]    io_imemAxi_ar_payload_prot,
  output wire          io_imemAxi_r_valid,
  input  wire          io_imemAxi_r_ready,
  output wire [31:0]   io_imemAxi_r_payload_data,
  output wire [1:0]    io_imemAxi_r_payload_resp,
  input  wire          io_dmemAxi_aw_valid,
  output wire          io_dmemAxi_aw_ready,
  input  wire [31:0]   io_dmemAxi_aw_payload_addr,
  input  wire [3:0]    io_dmemAxi_aw_payload_id,
  input  wire [7:0]    io_dmemAxi_aw_payload_len,
  input  wire [2:0]    io_dmemAxi_aw_payload_size,
  input  wire [1:0]    io_dmemAxi_aw_payload_burst,
  input  wire          io_dmemAxi_w_valid,
  output wire          io_dmemAxi_w_ready,
  input  wire [31:0]   io_dmemAxi_w_payload_data,
  input  wire [3:0]    io_dmemAxi_w_payload_strb,
  input  wire          io_dmemAxi_w_payload_last,
  output wire          io_dmemAxi_b_valid,
  input  wire          io_dmemAxi_b_ready,
  output wire [3:0]    io_dmemAxi_b_payload_id,
  output wire [1:0]    io_dmemAxi_b_payload_resp,
  input  wire          io_dmemAxi_ar_valid,
  output wire          io_dmemAxi_ar_ready,
  input  wire [31:0]   io_dmemAxi_ar_payload_addr,
  input  wire [3:0]    io_dmemAxi_ar_payload_id,
  input  wire [7:0]    io_dmemAxi_ar_payload_len,
  input  wire [2:0]    io_dmemAxi_ar_payload_size,
  input  wire [1:0]    io_dmemAxi_ar_payload_burst,
  output wire          io_dmemAxi_r_valid,
  input  wire          io_dmemAxi_r_ready,
  output wire [31:0]   io_dmemAxi_r_payload_data,
  output wire [3:0]    io_dmemAxi_r_payload_id,
  output wire [1:0]    io_dmemAxi_r_payload_resp,
  output wire          io_dmemAxi_r_payload_last,
  output wire          io_irq,
  input  wire          clk,
  input  wire          reset
);

  wire                cores_0_io_imemWrite_valid;
  wire                cores_0_io_dmemAxi_ar_valid;
  wire       [31:0]   cores_0_io_dmemAxi_ar_payload_addr;
  wire       [3:0]    cores_0_io_dmemAxi_ar_payload_id;
  wire       [7:0]    cores_0_io_dmemAxi_ar_payload_len;
  wire       [2:0]    cores_0_io_dmemAxi_ar_payload_size;
  wire       [1:0]    cores_0_io_dmemAxi_ar_payload_burst;
  wire                cores_0_io_dmemAxi_aw_valid;
  wire       [31:0]   cores_0_io_dmemAxi_aw_payload_addr;
  wire       [3:0]    cores_0_io_dmemAxi_aw_payload_id;
  wire       [7:0]    cores_0_io_dmemAxi_aw_payload_len;
  wire       [2:0]    cores_0_io_dmemAxi_aw_payload_size;
  wire       [1:0]    cores_0_io_dmemAxi_aw_payload_burst;
  wire                cores_0_io_dmemAxi_w_valid;
  wire       [31:0]   cores_0_io_dmemAxi_w_payload_data;
  wire       [3:0]    cores_0_io_dmemAxi_w_payload_strb;
  wire                cores_0_io_dmemAxi_w_payload_last;
  wire                cores_0_io_dmemAxi_r_ready;
  wire                cores_0_io_dmemAxi_b_ready;
  wire                cores_0_io_halted;
  wire                cores_0_io_running;
  wire       [9:0]    cores_0_io_pc;
  wire                cores_0_io_wawConflict;
  wire       [31:0]   cores_0_io_cycleCount;
  wire                memSub_io_corePorts_0_ar_ready;
  wire                memSub_io_corePorts_0_aw_ready;
  wire                memSub_io_corePorts_0_w_ready;
  wire                memSub_io_corePorts_0_r_valid;
  wire       [31:0]   memSub_io_corePorts_0_r_payload_data;
  wire       [3:0]    memSub_io_corePorts_0_r_payload_id;
  wire       [1:0]    memSub_io_corePorts_0_r_payload_resp;
  wire                memSub_io_corePorts_0_r_payload_last;
  wire                memSub_io_corePorts_0_b_valid;
  wire       [3:0]    memSub_io_corePorts_0_b_payload_id;
  wire       [1:0]    memSub_io_corePorts_0_b_payload_resp;
  wire                memSub_io_hostPort_ar_ready;
  wire                memSub_io_hostPort_aw_ready;
  wire                memSub_io_hostPort_w_ready;
  wire                memSub_io_hostPort_r_valid;
  wire       [31:0]   memSub_io_hostPort_r_payload_data;
  wire       [3:0]    memSub_io_hostPort_r_payload_id;
  wire       [1:0]    memSub_io_hostPort_r_payload_resp;
  wire                memSub_io_hostPort_r_payload_last;
  wire                memSub_io_hostPort_b_valid;
  wire       [3:0]    memSub_io_hostPort_b_payload_id;
  wire       [1:0]    memSub_io_hostPort_b_payload_resp;
  wire                hostIf_io_axiLite_aw_ready;
  wire                hostIf_io_axiLite_w_ready;
  wire                hostIf_io_axiLite_b_valid;
  wire       [1:0]    hostIf_io_axiLite_b_payload_resp;
  wire                hostIf_io_axiLite_ar_ready;
  wire                hostIf_io_axiLite_r_valid;
  wire       [31:0]   hostIf_io_axiLite_r_payload_data;
  wire       [1:0]    hostIf_io_axiLite_r_payload_resp;
  wire                hostIf_io_coreStart_0;
  wire                hostIf_io_coreReset_0;
  wire                hostIf_io_irq;
  wire       [29:0]   _zz_imemBusCtrl_wordIdx;
  wire       [26:0]   _zz_imemBusCtrl_instrAddr;
  wire       [7:0]    _zz_imemBusCtrl_accumulator_1;
  wire       [7:0]    _zz_imemBusCtrl_accumulator_2;
  wire       [7:0]    _zz_imemBusCtrl_accumulator_3;
  wire       [7:0]    _zz_imemBusCtrl_accumulator_4;
  wire       [7:0]    _zz_imemBusCtrl_accumulator_5;
  wire       [7:0]    _zz_imemBusCtrl_accumulator_6;
  wire       [7:0]    _zz_imemBusCtrl_accumulator_7;
  wire       [7:0]    _zz_imemBusCtrl_accumulator_8;
  wire       [7:0]    _zz_imemBusCtrl_accumulator_9;
  wire       [7:0]    _zz_imemBusCtrl_accumulator_10;
  wire       [7:0]    _zz_imemBusCtrl_accumulator_11;
  wire       [7:0]    _zz_imemBusCtrl_accumulator_12;
  wire       [7:0]    _zz_imemBusCtrl_accumulator_13;
  wire       [7:0]    _zz_imemBusCtrl_accumulator_14;
  wire       [7:0]    _zz_imemBusCtrl_accumulator_15;
  wire       [7:0]    _zz_imemBusCtrl_accumulator_16;
  wire       [7:0]    _zz_imemBusCtrl_accumulator_17;
  wire       [7:0]    _zz_imemBusCtrl_accumulator_18;
  wire       [7:0]    _zz_imemBusCtrl_accumulator_19;
  wire       [7:0]    _zz_imemBusCtrl_accumulator_20;
  wire       [7:0]    _zz_imemBusCtrl_accumulator_21;
  wire       [7:0]    _zz_imemBusCtrl_accumulator_22;
  wire       [7:0]    _zz_imemBusCtrl_accumulator_23;
  wire       [7:0]    _zz_imemBusCtrl_accumulator_24;
  wire       [7:0]    _zz_imemBusCtrl_accumulator_25;
  wire       [7:0]    _zz_imemBusCtrl_accumulator_26;
  wire       [7:0]    _zz_imemBusCtrl_accumulator_27;
  wire       [7:0]    _zz_imemBusCtrl_accumulator_28;
  wire       [7:0]    _zz_imemBusCtrl_accumulator_29;
  wire       [7:0]    _zz_imemBusCtrl_accumulator_30;
  wire       [7:0]    _zz_imemBusCtrl_accumulator_31;
  wire       [7:0]    _zz_imemBusCtrl_accumulator_32;
  wire       [7:0]    _zz_imemBusCtrl_accumulator_33;
  wire       [7:0]    _zz_imemBusCtrl_accumulator_34;
  wire       [7:0]    _zz_imemBusCtrl_accumulator_35;
  wire       [7:0]    _zz_imemBusCtrl_accumulator_36;
  wire       [7:0]    _zz_imemBusCtrl_accumulator_37;
  wire       [7:0]    _zz_imemBusCtrl_accumulator_38;
  wire       [7:0]    _zz_imemBusCtrl_accumulator_39;
  wire       [7:0]    _zz_imemBusCtrl_accumulator_40;
  wire       [7:0]    _zz_imemBusCtrl_accumulator_41;
  wire       [7:0]    _zz_imemBusCtrl_accumulator_42;
  wire       [7:0]    _zz_imemBusCtrl_accumulator_43;
  wire       [7:0]    _zz_imemBusCtrl_accumulator_44;
  wire       [7:0]    _zz_imemBusCtrl_accumulator_45;
  wire       [7:0]    _zz_imemBusCtrl_accumulator_46;
  wire       [7:0]    _zz_imemBusCtrl_accumulator_47;
  wire       [7:0]    _zz_imemBusCtrl_accumulator_48;
  wire       [7:0]    _zz_imemBusCtrl_accumulator_49;
  wire       [7:0]    _zz_imemBusCtrl_accumulator_50;
  wire       [7:0]    _zz_imemBusCtrl_accumulator_51;
  wire       [7:0]    _zz_imemBusCtrl_accumulator_52;
  wire       [7:0]    _zz_imemBusCtrl_accumulator_53;
  wire       [7:0]    _zz_imemBusCtrl_accumulator_54;
  wire       [7:0]    _zz_imemBusCtrl_accumulator_55;
  wire       [7:0]    _zz_imemBusCtrl_accumulator_56;
  wire       [7:0]    _zz_imemBusCtrl_accumulator_57;
  wire       [7:0]    _zz_imemBusCtrl_accumulator_58;
  wire       [7:0]    _zz_imemBusCtrl_accumulator_59;
  wire       [7:0]    _zz_imemBusCtrl_accumulator_60;
  wire       [7:0]    _zz_imemBusCtrl_accumulator_61;
  wire       [7:0]    _zz_imemBusCtrl_accumulator_62;
  wire       [7:0]    _zz_imemBusCtrl_accumulator_63;
  wire       [7:0]    _zz_imemBusCtrl_accumulator_64;
  wire       [7:0]    _zz_imemBusCtrl_commitData_1;
  wire       [7:0]    _zz_imemBusCtrl_commitData_2;
  wire       [7:0]    _zz_imemBusCtrl_commitData_3;
  wire       [7:0]    _zz_imemBusCtrl_commitData_4;
  wire       [7:0]    _zz_imemBusCtrl_commitData_5;
  wire       [7:0]    _zz_imemBusCtrl_commitData_6;
  wire       [7:0]    _zz_imemBusCtrl_commitData_7;
  wire       [7:0]    _zz_imemBusCtrl_commitData_8;
  wire       [7:0]    _zz_imemBusCtrl_commitData_9;
  wire       [7:0]    _zz_imemBusCtrl_commitData_10;
  wire       [7:0]    _zz_imemBusCtrl_commitData_11;
  wire       [7:0]    _zz_imemBusCtrl_commitData_12;
  wire       [7:0]    _zz_imemBusCtrl_commitData_13;
  wire       [7:0]    _zz_imemBusCtrl_commitData_14;
  wire       [7:0]    _zz_imemBusCtrl_commitData_15;
  wire       [7:0]    _zz_imemBusCtrl_commitData_16;
  wire       [7:0]    _zz_imemBusCtrl_commitData_17;
  wire       [7:0]    _zz_imemBusCtrl_commitData_18;
  wire       [7:0]    _zz_imemBusCtrl_commitData_19;
  wire       [7:0]    _zz_imemBusCtrl_commitData_20;
  wire       [7:0]    _zz_imemBusCtrl_commitData_21;
  wire       [7:0]    _zz_imemBusCtrl_commitData_22;
  wire       [7:0]    _zz_imemBusCtrl_commitData_23;
  wire       [7:0]    _zz_imemBusCtrl_commitData_24;
  wire       [7:0]    _zz_imemBusCtrl_commitData_25;
  wire       [7:0]    _zz_imemBusCtrl_commitData_26;
  wire       [7:0]    _zz_imemBusCtrl_commitData_27;
  wire       [7:0]    _zz_imemBusCtrl_commitData_28;
  wire       [7:0]    _zz_imemBusCtrl_commitData_29;
  wire       [7:0]    _zz_imemBusCtrl_commitData_30;
  wire       [7:0]    _zz_imemBusCtrl_commitData_31;
  wire       [7:0]    _zz_imemBusCtrl_commitData_32;
  wire       [7:0]    _zz_imemBusCtrl_commitData_33;
  wire       [7:0]    _zz_imemBusCtrl_commitData_34;
  wire       [7:0]    _zz_imemBusCtrl_commitData_35;
  wire       [7:0]    _zz_imemBusCtrl_commitData_36;
  wire       [7:0]    _zz_imemBusCtrl_commitData_37;
  wire       [7:0]    _zz_imemBusCtrl_commitData_38;
  wire       [7:0]    _zz_imemBusCtrl_commitData_39;
  wire       [7:0]    _zz_imemBusCtrl_commitData_40;
  wire       [7:0]    _zz_imemBusCtrl_commitData_41;
  wire       [7:0]    _zz_imemBusCtrl_commitData_42;
  wire       [7:0]    _zz_imemBusCtrl_commitData_43;
  wire       [7:0]    _zz_imemBusCtrl_commitData_44;
  wire       [7:0]    _zz_imemBusCtrl_commitData_45;
  wire       [7:0]    _zz_imemBusCtrl_commitData_46;
  wire       [7:0]    _zz_imemBusCtrl_commitData_47;
  wire       [7:0]    _zz_imemBusCtrl_commitData_48;
  wire       [7:0]    _zz_imemBusCtrl_commitData_49;
  wire       [7:0]    _zz_imemBusCtrl_commitData_50;
  wire       [7:0]    _zz_imemBusCtrl_commitData_51;
  wire       [7:0]    _zz_imemBusCtrl_commitData_52;
  wire       [7:0]    _zz_imemBusCtrl_commitData_53;
  wire       [7:0]    _zz_imemBusCtrl_commitData_54;
  wire       [7:0]    _zz_imemBusCtrl_commitData_55;
  wire       [7:0]    _zz_imemBusCtrl_commitData_56;
  wire       [7:0]    _zz_imemBusCtrl_commitData_57;
  wire       [7:0]    _zz_imemBusCtrl_commitData_58;
  wire       [7:0]    _zz_imemBusCtrl_commitData_59;
  wire       [7:0]    _zz_imemBusCtrl_commitData_60;
  wire       [7:0]    _zz_imemBusCtrl_commitData_61;
  wire       [7:0]    _zz_imemBusCtrl_commitData_62;
  wire       [7:0]    _zz_imemBusCtrl_commitData_63;
  wire       [7:0]    _zz_imemBusCtrl_commitData_64;
  reg                 imemBusCtrl_awReady;
  reg                 imemBusCtrl_wReady;
  reg                 imemBusCtrl_bValid;
  reg        [31:0]   imemBusCtrl_awAddr;
  reg        [31:0]   imemBusCtrl_wData;
  wire                imemBusCtrl_awFire;
  wire                imemBusCtrl_wFire;
  reg                 imemBusCtrl_bothFired;
  reg                 imemBusCtrl_awDone;
  reg                 imemBusCtrl_wDone;
  wire                when_VliwSimdSoc_l135;
  wire                when_VliwSimdSoc_l149;
  wire                when_VliwSimdSoc_l156;
  reg        [255:0]  imemBusCtrl_accumulator;
  wire       [2:0]    imemBusCtrl_wordIdx;
  wire       [9:0]    imemBusCtrl_instrAddr;
  wire       [0:0]    imemBusCtrl_coreSelect;
  wire                imemBusCtrl_isLastWord;
  wire       [8:0]    _zz_imemBusCtrl_accumulator;
  reg                 imemBusCtrl_commitValid;
  reg        [9:0]    imemBusCtrl_commitAddr;
  reg        [0:0]    imemBusCtrl_commitCore;
  reg        [255:0]  imemBusCtrl_commitData;
  wire                when_VliwSimdSoc_l204;
  wire       [8:0]    _zz_imemBusCtrl_commitData;
  wire                when_VliwSimdSoc_l228;

  assign _zz_imemBusCtrl_wordIdx = (imemBusCtrl_awAddr >>> 2'd2);
  assign _zz_imemBusCtrl_instrAddr = (imemBusCtrl_awAddr >>> 3'd5);
  assign _zz_imemBusCtrl_accumulator_1 = (_zz_imemBusCtrl_accumulator_2 + 8'h0);
  assign _zz_imemBusCtrl_accumulator_2 = _zz_imemBusCtrl_accumulator[7:0];
  assign _zz_imemBusCtrl_accumulator_3 = (_zz_imemBusCtrl_accumulator_4 + 8'h01);
  assign _zz_imemBusCtrl_accumulator_4 = _zz_imemBusCtrl_accumulator[7:0];
  assign _zz_imemBusCtrl_accumulator_5 = (_zz_imemBusCtrl_accumulator_6 + 8'h02);
  assign _zz_imemBusCtrl_accumulator_6 = _zz_imemBusCtrl_accumulator[7:0];
  assign _zz_imemBusCtrl_accumulator_7 = (_zz_imemBusCtrl_accumulator_8 + 8'h03);
  assign _zz_imemBusCtrl_accumulator_8 = _zz_imemBusCtrl_accumulator[7:0];
  assign _zz_imemBusCtrl_accumulator_9 = (_zz_imemBusCtrl_accumulator_10 + 8'h04);
  assign _zz_imemBusCtrl_accumulator_10 = _zz_imemBusCtrl_accumulator[7:0];
  assign _zz_imemBusCtrl_accumulator_11 = (_zz_imemBusCtrl_accumulator_12 + 8'h05);
  assign _zz_imemBusCtrl_accumulator_12 = _zz_imemBusCtrl_accumulator[7:0];
  assign _zz_imemBusCtrl_accumulator_13 = (_zz_imemBusCtrl_accumulator_14 + 8'h06);
  assign _zz_imemBusCtrl_accumulator_14 = _zz_imemBusCtrl_accumulator[7:0];
  assign _zz_imemBusCtrl_accumulator_15 = (_zz_imemBusCtrl_accumulator_16 + 8'h07);
  assign _zz_imemBusCtrl_accumulator_16 = _zz_imemBusCtrl_accumulator[7:0];
  assign _zz_imemBusCtrl_accumulator_17 = (_zz_imemBusCtrl_accumulator_18 + 8'h08);
  assign _zz_imemBusCtrl_accumulator_18 = _zz_imemBusCtrl_accumulator[7:0];
  assign _zz_imemBusCtrl_accumulator_19 = (_zz_imemBusCtrl_accumulator_20 + 8'h09);
  assign _zz_imemBusCtrl_accumulator_20 = _zz_imemBusCtrl_accumulator[7:0];
  assign _zz_imemBusCtrl_accumulator_21 = (_zz_imemBusCtrl_accumulator_22 + 8'h0a);
  assign _zz_imemBusCtrl_accumulator_22 = _zz_imemBusCtrl_accumulator[7:0];
  assign _zz_imemBusCtrl_accumulator_23 = (_zz_imemBusCtrl_accumulator_24 + 8'h0b);
  assign _zz_imemBusCtrl_accumulator_24 = _zz_imemBusCtrl_accumulator[7:0];
  assign _zz_imemBusCtrl_accumulator_25 = (_zz_imemBusCtrl_accumulator_26 + 8'h0c);
  assign _zz_imemBusCtrl_accumulator_26 = _zz_imemBusCtrl_accumulator[7:0];
  assign _zz_imemBusCtrl_accumulator_27 = (_zz_imemBusCtrl_accumulator_28 + 8'h0d);
  assign _zz_imemBusCtrl_accumulator_28 = _zz_imemBusCtrl_accumulator[7:0];
  assign _zz_imemBusCtrl_accumulator_29 = (_zz_imemBusCtrl_accumulator_30 + 8'h0e);
  assign _zz_imemBusCtrl_accumulator_30 = _zz_imemBusCtrl_accumulator[7:0];
  assign _zz_imemBusCtrl_accumulator_31 = (_zz_imemBusCtrl_accumulator_32 + 8'h0f);
  assign _zz_imemBusCtrl_accumulator_32 = _zz_imemBusCtrl_accumulator[7:0];
  assign _zz_imemBusCtrl_accumulator_33 = (_zz_imemBusCtrl_accumulator_34 + 8'h10);
  assign _zz_imemBusCtrl_accumulator_34 = _zz_imemBusCtrl_accumulator[7:0];
  assign _zz_imemBusCtrl_accumulator_35 = (_zz_imemBusCtrl_accumulator_36 + 8'h11);
  assign _zz_imemBusCtrl_accumulator_36 = _zz_imemBusCtrl_accumulator[7:0];
  assign _zz_imemBusCtrl_accumulator_37 = (_zz_imemBusCtrl_accumulator_38 + 8'h12);
  assign _zz_imemBusCtrl_accumulator_38 = _zz_imemBusCtrl_accumulator[7:0];
  assign _zz_imemBusCtrl_accumulator_39 = (_zz_imemBusCtrl_accumulator_40 + 8'h13);
  assign _zz_imemBusCtrl_accumulator_40 = _zz_imemBusCtrl_accumulator[7:0];
  assign _zz_imemBusCtrl_accumulator_41 = (_zz_imemBusCtrl_accumulator_42 + 8'h14);
  assign _zz_imemBusCtrl_accumulator_42 = _zz_imemBusCtrl_accumulator[7:0];
  assign _zz_imemBusCtrl_accumulator_43 = (_zz_imemBusCtrl_accumulator_44 + 8'h15);
  assign _zz_imemBusCtrl_accumulator_44 = _zz_imemBusCtrl_accumulator[7:0];
  assign _zz_imemBusCtrl_accumulator_45 = (_zz_imemBusCtrl_accumulator_46 + 8'h16);
  assign _zz_imemBusCtrl_accumulator_46 = _zz_imemBusCtrl_accumulator[7:0];
  assign _zz_imemBusCtrl_accumulator_47 = (_zz_imemBusCtrl_accumulator_48 + 8'h17);
  assign _zz_imemBusCtrl_accumulator_48 = _zz_imemBusCtrl_accumulator[7:0];
  assign _zz_imemBusCtrl_accumulator_49 = (_zz_imemBusCtrl_accumulator_50 + 8'h18);
  assign _zz_imemBusCtrl_accumulator_50 = _zz_imemBusCtrl_accumulator[7:0];
  assign _zz_imemBusCtrl_accumulator_51 = (_zz_imemBusCtrl_accumulator_52 + 8'h19);
  assign _zz_imemBusCtrl_accumulator_52 = _zz_imemBusCtrl_accumulator[7:0];
  assign _zz_imemBusCtrl_accumulator_53 = (_zz_imemBusCtrl_accumulator_54 + 8'h1a);
  assign _zz_imemBusCtrl_accumulator_54 = _zz_imemBusCtrl_accumulator[7:0];
  assign _zz_imemBusCtrl_accumulator_55 = (_zz_imemBusCtrl_accumulator_56 + 8'h1b);
  assign _zz_imemBusCtrl_accumulator_56 = _zz_imemBusCtrl_accumulator[7:0];
  assign _zz_imemBusCtrl_accumulator_57 = (_zz_imemBusCtrl_accumulator_58 + 8'h1c);
  assign _zz_imemBusCtrl_accumulator_58 = _zz_imemBusCtrl_accumulator[7:0];
  assign _zz_imemBusCtrl_accumulator_59 = (_zz_imemBusCtrl_accumulator_60 + 8'h1d);
  assign _zz_imemBusCtrl_accumulator_60 = _zz_imemBusCtrl_accumulator[7:0];
  assign _zz_imemBusCtrl_accumulator_61 = (_zz_imemBusCtrl_accumulator_62 + 8'h1e);
  assign _zz_imemBusCtrl_accumulator_62 = _zz_imemBusCtrl_accumulator[7:0];
  assign _zz_imemBusCtrl_accumulator_63 = (_zz_imemBusCtrl_accumulator_64 + 8'h1f);
  assign _zz_imemBusCtrl_accumulator_64 = _zz_imemBusCtrl_accumulator[7:0];
  assign _zz_imemBusCtrl_commitData_1 = (_zz_imemBusCtrl_commitData_2 + 8'h0);
  assign _zz_imemBusCtrl_commitData_2 = _zz_imemBusCtrl_commitData[7:0];
  assign _zz_imemBusCtrl_commitData_3 = (_zz_imemBusCtrl_commitData_4 + 8'h01);
  assign _zz_imemBusCtrl_commitData_4 = _zz_imemBusCtrl_commitData[7:0];
  assign _zz_imemBusCtrl_commitData_5 = (_zz_imemBusCtrl_commitData_6 + 8'h02);
  assign _zz_imemBusCtrl_commitData_6 = _zz_imemBusCtrl_commitData[7:0];
  assign _zz_imemBusCtrl_commitData_7 = (_zz_imemBusCtrl_commitData_8 + 8'h03);
  assign _zz_imemBusCtrl_commitData_8 = _zz_imemBusCtrl_commitData[7:0];
  assign _zz_imemBusCtrl_commitData_9 = (_zz_imemBusCtrl_commitData_10 + 8'h04);
  assign _zz_imemBusCtrl_commitData_10 = _zz_imemBusCtrl_commitData[7:0];
  assign _zz_imemBusCtrl_commitData_11 = (_zz_imemBusCtrl_commitData_12 + 8'h05);
  assign _zz_imemBusCtrl_commitData_12 = _zz_imemBusCtrl_commitData[7:0];
  assign _zz_imemBusCtrl_commitData_13 = (_zz_imemBusCtrl_commitData_14 + 8'h06);
  assign _zz_imemBusCtrl_commitData_14 = _zz_imemBusCtrl_commitData[7:0];
  assign _zz_imemBusCtrl_commitData_15 = (_zz_imemBusCtrl_commitData_16 + 8'h07);
  assign _zz_imemBusCtrl_commitData_16 = _zz_imemBusCtrl_commitData[7:0];
  assign _zz_imemBusCtrl_commitData_17 = (_zz_imemBusCtrl_commitData_18 + 8'h08);
  assign _zz_imemBusCtrl_commitData_18 = _zz_imemBusCtrl_commitData[7:0];
  assign _zz_imemBusCtrl_commitData_19 = (_zz_imemBusCtrl_commitData_20 + 8'h09);
  assign _zz_imemBusCtrl_commitData_20 = _zz_imemBusCtrl_commitData[7:0];
  assign _zz_imemBusCtrl_commitData_21 = (_zz_imemBusCtrl_commitData_22 + 8'h0a);
  assign _zz_imemBusCtrl_commitData_22 = _zz_imemBusCtrl_commitData[7:0];
  assign _zz_imemBusCtrl_commitData_23 = (_zz_imemBusCtrl_commitData_24 + 8'h0b);
  assign _zz_imemBusCtrl_commitData_24 = _zz_imemBusCtrl_commitData[7:0];
  assign _zz_imemBusCtrl_commitData_25 = (_zz_imemBusCtrl_commitData_26 + 8'h0c);
  assign _zz_imemBusCtrl_commitData_26 = _zz_imemBusCtrl_commitData[7:0];
  assign _zz_imemBusCtrl_commitData_27 = (_zz_imemBusCtrl_commitData_28 + 8'h0d);
  assign _zz_imemBusCtrl_commitData_28 = _zz_imemBusCtrl_commitData[7:0];
  assign _zz_imemBusCtrl_commitData_29 = (_zz_imemBusCtrl_commitData_30 + 8'h0e);
  assign _zz_imemBusCtrl_commitData_30 = _zz_imemBusCtrl_commitData[7:0];
  assign _zz_imemBusCtrl_commitData_31 = (_zz_imemBusCtrl_commitData_32 + 8'h0f);
  assign _zz_imemBusCtrl_commitData_32 = _zz_imemBusCtrl_commitData[7:0];
  assign _zz_imemBusCtrl_commitData_33 = (_zz_imemBusCtrl_commitData_34 + 8'h10);
  assign _zz_imemBusCtrl_commitData_34 = _zz_imemBusCtrl_commitData[7:0];
  assign _zz_imemBusCtrl_commitData_35 = (_zz_imemBusCtrl_commitData_36 + 8'h11);
  assign _zz_imemBusCtrl_commitData_36 = _zz_imemBusCtrl_commitData[7:0];
  assign _zz_imemBusCtrl_commitData_37 = (_zz_imemBusCtrl_commitData_38 + 8'h12);
  assign _zz_imemBusCtrl_commitData_38 = _zz_imemBusCtrl_commitData[7:0];
  assign _zz_imemBusCtrl_commitData_39 = (_zz_imemBusCtrl_commitData_40 + 8'h13);
  assign _zz_imemBusCtrl_commitData_40 = _zz_imemBusCtrl_commitData[7:0];
  assign _zz_imemBusCtrl_commitData_41 = (_zz_imemBusCtrl_commitData_42 + 8'h14);
  assign _zz_imemBusCtrl_commitData_42 = _zz_imemBusCtrl_commitData[7:0];
  assign _zz_imemBusCtrl_commitData_43 = (_zz_imemBusCtrl_commitData_44 + 8'h15);
  assign _zz_imemBusCtrl_commitData_44 = _zz_imemBusCtrl_commitData[7:0];
  assign _zz_imemBusCtrl_commitData_45 = (_zz_imemBusCtrl_commitData_46 + 8'h16);
  assign _zz_imemBusCtrl_commitData_46 = _zz_imemBusCtrl_commitData[7:0];
  assign _zz_imemBusCtrl_commitData_47 = (_zz_imemBusCtrl_commitData_48 + 8'h17);
  assign _zz_imemBusCtrl_commitData_48 = _zz_imemBusCtrl_commitData[7:0];
  assign _zz_imemBusCtrl_commitData_49 = (_zz_imemBusCtrl_commitData_50 + 8'h18);
  assign _zz_imemBusCtrl_commitData_50 = _zz_imemBusCtrl_commitData[7:0];
  assign _zz_imemBusCtrl_commitData_51 = (_zz_imemBusCtrl_commitData_52 + 8'h19);
  assign _zz_imemBusCtrl_commitData_52 = _zz_imemBusCtrl_commitData[7:0];
  assign _zz_imemBusCtrl_commitData_53 = (_zz_imemBusCtrl_commitData_54 + 8'h1a);
  assign _zz_imemBusCtrl_commitData_54 = _zz_imemBusCtrl_commitData[7:0];
  assign _zz_imemBusCtrl_commitData_55 = (_zz_imemBusCtrl_commitData_56 + 8'h1b);
  assign _zz_imemBusCtrl_commitData_56 = _zz_imemBusCtrl_commitData[7:0];
  assign _zz_imemBusCtrl_commitData_57 = (_zz_imemBusCtrl_commitData_58 + 8'h1c);
  assign _zz_imemBusCtrl_commitData_58 = _zz_imemBusCtrl_commitData[7:0];
  assign _zz_imemBusCtrl_commitData_59 = (_zz_imemBusCtrl_commitData_60 + 8'h1d);
  assign _zz_imemBusCtrl_commitData_60 = _zz_imemBusCtrl_commitData[7:0];
  assign _zz_imemBusCtrl_commitData_61 = (_zz_imemBusCtrl_commitData_62 + 8'h1e);
  assign _zz_imemBusCtrl_commitData_62 = _zz_imemBusCtrl_commitData[7:0];
  assign _zz_imemBusCtrl_commitData_63 = (_zz_imemBusCtrl_commitData_64 + 8'h1f);
  assign _zz_imemBusCtrl_commitData_64 = _zz_imemBusCtrl_commitData[7:0];
  VliwCore cores_0 (
    .io_imemWrite_valid          (cores_0_io_imemWrite_valid                ), //i
    .io_imemWrite_payload_addr   (imemBusCtrl_commitAddr[9:0]               ), //i
    .io_imemWrite_payload_data   (imemBusCtrl_commitData[255:0]             ), //i
    .io_dmemAxi_aw_valid         (cores_0_io_dmemAxi_aw_valid               ), //o
    .io_dmemAxi_aw_ready         (memSub_io_corePorts_0_aw_ready            ), //i
    .io_dmemAxi_aw_payload_addr  (cores_0_io_dmemAxi_aw_payload_addr[31:0]  ), //o
    .io_dmemAxi_aw_payload_id    (cores_0_io_dmemAxi_aw_payload_id[3:0]     ), //o
    .io_dmemAxi_aw_payload_len   (cores_0_io_dmemAxi_aw_payload_len[7:0]    ), //o
    .io_dmemAxi_aw_payload_size  (cores_0_io_dmemAxi_aw_payload_size[2:0]   ), //o
    .io_dmemAxi_aw_payload_burst (cores_0_io_dmemAxi_aw_payload_burst[1:0]  ), //o
    .io_dmemAxi_w_valid          (cores_0_io_dmemAxi_w_valid                ), //o
    .io_dmemAxi_w_ready          (memSub_io_corePorts_0_w_ready             ), //i
    .io_dmemAxi_w_payload_data   (cores_0_io_dmemAxi_w_payload_data[31:0]   ), //o
    .io_dmemAxi_w_payload_strb   (cores_0_io_dmemAxi_w_payload_strb[3:0]    ), //o
    .io_dmemAxi_w_payload_last   (cores_0_io_dmemAxi_w_payload_last         ), //o
    .io_dmemAxi_b_valid          (memSub_io_corePorts_0_b_valid             ), //i
    .io_dmemAxi_b_ready          (cores_0_io_dmemAxi_b_ready                ), //o
    .io_dmemAxi_b_payload_id     (memSub_io_corePorts_0_b_payload_id[3:0]   ), //i
    .io_dmemAxi_b_payload_resp   (memSub_io_corePorts_0_b_payload_resp[1:0] ), //i
    .io_dmemAxi_ar_valid         (cores_0_io_dmemAxi_ar_valid               ), //o
    .io_dmemAxi_ar_ready         (memSub_io_corePorts_0_ar_ready            ), //i
    .io_dmemAxi_ar_payload_addr  (cores_0_io_dmemAxi_ar_payload_addr[31:0]  ), //o
    .io_dmemAxi_ar_payload_id    (cores_0_io_dmemAxi_ar_payload_id[3:0]     ), //o
    .io_dmemAxi_ar_payload_len   (cores_0_io_dmemAxi_ar_payload_len[7:0]    ), //o
    .io_dmemAxi_ar_payload_size  (cores_0_io_dmemAxi_ar_payload_size[2:0]   ), //o
    .io_dmemAxi_ar_payload_burst (cores_0_io_dmemAxi_ar_payload_burst[1:0]  ), //o
    .io_dmemAxi_r_valid          (memSub_io_corePorts_0_r_valid             ), //i
    .io_dmemAxi_r_ready          (cores_0_io_dmemAxi_r_ready                ), //o
    .io_dmemAxi_r_payload_data   (memSub_io_corePorts_0_r_payload_data[31:0]), //i
    .io_dmemAxi_r_payload_id     (memSub_io_corePorts_0_r_payload_id[3:0]   ), //i
    .io_dmemAxi_r_payload_resp   (memSub_io_corePorts_0_r_payload_resp[1:0] ), //i
    .io_dmemAxi_r_payload_last   (memSub_io_corePorts_0_r_payload_last      ), //i
    .io_start                    (hostIf_io_coreStart_0                     ), //i
    .io_halted                   (cores_0_io_halted                         ), //o
    .io_running                  (cores_0_io_running                        ), //o
    .io_pc                       (cores_0_io_pc[9:0]                        ), //o
    .io_wawConflict              (cores_0_io_wawConflict                    ), //o
    .io_cycleCount               (cores_0_io_cycleCount[31:0]               ), //o
    .clk                         (clk                                       ), //i
    .reset                       (reset                                     )  //i
  );
  MemorySubsystem memSub (
    .io_corePorts_0_aw_valid         (cores_0_io_dmemAxi_aw_valid               ), //i
    .io_corePorts_0_aw_ready         (memSub_io_corePorts_0_aw_ready            ), //o
    .io_corePorts_0_aw_payload_addr  (cores_0_io_dmemAxi_aw_payload_addr[31:0]  ), //i
    .io_corePorts_0_aw_payload_id    (cores_0_io_dmemAxi_aw_payload_id[3:0]     ), //i
    .io_corePorts_0_aw_payload_len   (cores_0_io_dmemAxi_aw_payload_len[7:0]    ), //i
    .io_corePorts_0_aw_payload_size  (cores_0_io_dmemAxi_aw_payload_size[2:0]   ), //i
    .io_corePorts_0_aw_payload_burst (cores_0_io_dmemAxi_aw_payload_burst[1:0]  ), //i
    .io_corePorts_0_w_valid          (cores_0_io_dmemAxi_w_valid                ), //i
    .io_corePorts_0_w_ready          (memSub_io_corePorts_0_w_ready             ), //o
    .io_corePorts_0_w_payload_data   (cores_0_io_dmemAxi_w_payload_data[31:0]   ), //i
    .io_corePorts_0_w_payload_strb   (cores_0_io_dmemAxi_w_payload_strb[3:0]    ), //i
    .io_corePorts_0_w_payload_last   (cores_0_io_dmemAxi_w_payload_last         ), //i
    .io_corePorts_0_b_valid          (memSub_io_corePorts_0_b_valid             ), //o
    .io_corePorts_0_b_ready          (cores_0_io_dmemAxi_b_ready                ), //i
    .io_corePorts_0_b_payload_id     (memSub_io_corePorts_0_b_payload_id[3:0]   ), //o
    .io_corePorts_0_b_payload_resp   (memSub_io_corePorts_0_b_payload_resp[1:0] ), //o
    .io_corePorts_0_ar_valid         (cores_0_io_dmemAxi_ar_valid               ), //i
    .io_corePorts_0_ar_ready         (memSub_io_corePorts_0_ar_ready            ), //o
    .io_corePorts_0_ar_payload_addr  (cores_0_io_dmemAxi_ar_payload_addr[31:0]  ), //i
    .io_corePorts_0_ar_payload_id    (cores_0_io_dmemAxi_ar_payload_id[3:0]     ), //i
    .io_corePorts_0_ar_payload_len   (cores_0_io_dmemAxi_ar_payload_len[7:0]    ), //i
    .io_corePorts_0_ar_payload_size  (cores_0_io_dmemAxi_ar_payload_size[2:0]   ), //i
    .io_corePorts_0_ar_payload_burst (cores_0_io_dmemAxi_ar_payload_burst[1:0]  ), //i
    .io_corePorts_0_r_valid          (memSub_io_corePorts_0_r_valid             ), //o
    .io_corePorts_0_r_ready          (cores_0_io_dmemAxi_r_ready                ), //i
    .io_corePorts_0_r_payload_data   (memSub_io_corePorts_0_r_payload_data[31:0]), //o
    .io_corePorts_0_r_payload_id     (memSub_io_corePorts_0_r_payload_id[3:0]   ), //o
    .io_corePorts_0_r_payload_resp   (memSub_io_corePorts_0_r_payload_resp[1:0] ), //o
    .io_corePorts_0_r_payload_last   (memSub_io_corePorts_0_r_payload_last      ), //o
    .io_hostPort_aw_valid            (io_dmemAxi_aw_valid                       ), //i
    .io_hostPort_aw_ready            (memSub_io_hostPort_aw_ready               ), //o
    .io_hostPort_aw_payload_addr     (io_dmemAxi_aw_payload_addr[31:0]          ), //i
    .io_hostPort_aw_payload_id       (io_dmemAxi_aw_payload_id[3:0]             ), //i
    .io_hostPort_aw_payload_len      (io_dmemAxi_aw_payload_len[7:0]            ), //i
    .io_hostPort_aw_payload_size     (io_dmemAxi_aw_payload_size[2:0]           ), //i
    .io_hostPort_aw_payload_burst    (io_dmemAxi_aw_payload_burst[1:0]          ), //i
    .io_hostPort_w_valid             (io_dmemAxi_w_valid                        ), //i
    .io_hostPort_w_ready             (memSub_io_hostPort_w_ready                ), //o
    .io_hostPort_w_payload_data      (io_dmemAxi_w_payload_data[31:0]           ), //i
    .io_hostPort_w_payload_strb      (io_dmemAxi_w_payload_strb[3:0]            ), //i
    .io_hostPort_w_payload_last      (io_dmemAxi_w_payload_last                 ), //i
    .io_hostPort_b_valid             (memSub_io_hostPort_b_valid                ), //o
    .io_hostPort_b_ready             (io_dmemAxi_b_ready                        ), //i
    .io_hostPort_b_payload_id        (memSub_io_hostPort_b_payload_id[3:0]      ), //o
    .io_hostPort_b_payload_resp      (memSub_io_hostPort_b_payload_resp[1:0]    ), //o
    .io_hostPort_ar_valid            (io_dmemAxi_ar_valid                       ), //i
    .io_hostPort_ar_ready            (memSub_io_hostPort_ar_ready               ), //o
    .io_hostPort_ar_payload_addr     (io_dmemAxi_ar_payload_addr[31:0]          ), //i
    .io_hostPort_ar_payload_id       (io_dmemAxi_ar_payload_id[3:0]             ), //i
    .io_hostPort_ar_payload_len      (io_dmemAxi_ar_payload_len[7:0]            ), //i
    .io_hostPort_ar_payload_size     (io_dmemAxi_ar_payload_size[2:0]           ), //i
    .io_hostPort_ar_payload_burst    (io_dmemAxi_ar_payload_burst[1:0]          ), //i
    .io_hostPort_r_valid             (memSub_io_hostPort_r_valid                ), //o
    .io_hostPort_r_ready             (io_dmemAxi_r_ready                        ), //i
    .io_hostPort_r_payload_data      (memSub_io_hostPort_r_payload_data[31:0]   ), //o
    .io_hostPort_r_payload_id        (memSub_io_hostPort_r_payload_id[3:0]      ), //o
    .io_hostPort_r_payload_resp      (memSub_io_hostPort_r_payload_resp[1:0]    ), //o
    .io_hostPort_r_payload_last      (memSub_io_hostPort_r_payload_last         ), //o
    .clk                             (clk                                       ), //i
    .reset                           (reset                                     )  //i
  );
  HostInterface hostIf (
    .io_axiLite_aw_valid        (io_csrAxi_aw_valid                    ), //i
    .io_axiLite_aw_ready        (hostIf_io_axiLite_aw_ready            ), //o
    .io_axiLite_aw_payload_addr (io_csrAxi_aw_payload_addr[31:0]       ), //i
    .io_axiLite_aw_payload_prot (io_csrAxi_aw_payload_prot[2:0]        ), //i
    .io_axiLite_w_valid         (io_csrAxi_w_valid                     ), //i
    .io_axiLite_w_ready         (hostIf_io_axiLite_w_ready             ), //o
    .io_axiLite_w_payload_data  (io_csrAxi_w_payload_data[31:0]        ), //i
    .io_axiLite_w_payload_strb  (io_csrAxi_w_payload_strb[3:0]         ), //i
    .io_axiLite_b_valid         (hostIf_io_axiLite_b_valid             ), //o
    .io_axiLite_b_ready         (io_csrAxi_b_ready                     ), //i
    .io_axiLite_b_payload_resp  (hostIf_io_axiLite_b_payload_resp[1:0] ), //o
    .io_axiLite_ar_valid        (io_csrAxi_ar_valid                    ), //i
    .io_axiLite_ar_ready        (hostIf_io_axiLite_ar_ready            ), //o
    .io_axiLite_ar_payload_addr (io_csrAxi_ar_payload_addr[31:0]       ), //i
    .io_axiLite_ar_payload_prot (io_csrAxi_ar_payload_prot[2:0]        ), //i
    .io_axiLite_r_valid         (hostIf_io_axiLite_r_valid             ), //o
    .io_axiLite_r_ready         (io_csrAxi_r_ready                     ), //i
    .io_axiLite_r_payload_data  (hostIf_io_axiLite_r_payload_data[31:0]), //o
    .io_axiLite_r_payload_resp  (hostIf_io_axiLite_r_payload_resp[1:0] ), //o
    .io_coreStart_0             (hostIf_io_coreStart_0                 ), //o
    .io_coreReset_0             (hostIf_io_coreReset_0                 ), //o
    .io_coreHalted_0            (cores_0_io_halted                     ), //i
    .io_coreRunning_0           (cores_0_io_running                    ), //i
    .io_corePc_0                (cores_0_io_pc[9:0]                    ), //i
    .io_coreCycles_0            (cores_0_io_cycleCount[31:0]           ), //i
    .io_irq                     (hostIf_io_irq                         ), //o
    .clk                        (clk                                   ), //i
    .reset                      (reset                                 )  //i
  );
  assign io_dmemAxi_aw_ready = memSub_io_hostPort_aw_ready;
  assign io_dmemAxi_w_ready = memSub_io_hostPort_w_ready;
  assign io_dmemAxi_b_valid = memSub_io_hostPort_b_valid;
  assign io_dmemAxi_b_payload_id = memSub_io_hostPort_b_payload_id;
  assign io_dmemAxi_b_payload_resp = memSub_io_hostPort_b_payload_resp;
  assign io_dmemAxi_ar_ready = memSub_io_hostPort_ar_ready;
  assign io_dmemAxi_r_valid = memSub_io_hostPort_r_valid;
  assign io_dmemAxi_r_payload_data = memSub_io_hostPort_r_payload_data;
  assign io_dmemAxi_r_payload_id = memSub_io_hostPort_r_payload_id;
  assign io_dmemAxi_r_payload_resp = memSub_io_hostPort_r_payload_resp;
  assign io_dmemAxi_r_payload_last = memSub_io_hostPort_r_payload_last;
  assign io_csrAxi_aw_ready = hostIf_io_axiLite_aw_ready;
  assign io_csrAxi_w_ready = hostIf_io_axiLite_w_ready;
  assign io_csrAxi_b_valid = hostIf_io_axiLite_b_valid;
  assign io_csrAxi_b_payload_resp = hostIf_io_axiLite_b_payload_resp;
  assign io_csrAxi_ar_ready = hostIf_io_axiLite_ar_ready;
  assign io_csrAxi_r_valid = hostIf_io_axiLite_r_valid;
  assign io_csrAxi_r_payload_data = hostIf_io_axiLite_r_payload_data;
  assign io_csrAxi_r_payload_resp = hostIf_io_axiLite_r_payload_resp;
  assign io_irq = hostIf_io_irq;
  assign io_imemAxi_aw_ready = imemBusCtrl_awReady;
  assign io_imemAxi_w_ready = imemBusCtrl_wReady;
  assign io_imemAxi_b_valid = imemBusCtrl_bValid;
  assign io_imemAxi_b_payload_resp = 2'b00;
  assign io_imemAxi_ar_ready = 1'b0;
  assign io_imemAxi_r_valid = 1'b0;
  assign io_imemAxi_r_payload_data = 32'h0;
  assign io_imemAxi_r_payload_resp = 2'b00;
  assign imemBusCtrl_awFire = (io_imemAxi_aw_valid && io_imemAxi_aw_ready);
  assign imemBusCtrl_wFire = (io_imemAxi_w_valid && io_imemAxi_w_ready);
  assign when_VliwSimdSoc_l135 = (imemBusCtrl_awFire && imemBusCtrl_wFire);
  assign when_VliwSimdSoc_l149 = (imemBusCtrl_awDone && imemBusCtrl_wFire);
  assign when_VliwSimdSoc_l156 = (imemBusCtrl_wDone && imemBusCtrl_awFire);
  assign imemBusCtrl_wordIdx = _zz_imemBusCtrl_wordIdx[2:0];
  assign imemBusCtrl_instrAddr = _zz_imemBusCtrl_instrAddr[9:0];
  assign imemBusCtrl_coreSelect = 1'b0;
  assign imemBusCtrl_isLastWord = (imemBusCtrl_wordIdx == 3'b111);
  assign _zz_imemBusCtrl_accumulator = (imemBusCtrl_wordIdx * 6'h20);
  assign when_VliwSimdSoc_l204 = (imemBusCtrl_bothFired && imemBusCtrl_isLastWord);
  assign _zz_imemBusCtrl_commitData = (imemBusCtrl_wordIdx * 6'h20);
  assign cores_0_io_imemWrite_valid = (imemBusCtrl_commitValid && 1'b1);
  assign when_VliwSimdSoc_l228 = (io_imemAxi_b_valid && io_imemAxi_b_ready);
  always @(posedge clk) begin
    if(reset) begin
      imemBusCtrl_awReady <= 1'b1;
      imemBusCtrl_wReady <= 1'b1;
      imemBusCtrl_bValid <= 1'b0;
      imemBusCtrl_bothFired <= 1'b0;
      imemBusCtrl_awDone <= 1'b0;
      imemBusCtrl_wDone <= 1'b0;
      imemBusCtrl_accumulator <= 256'h0;
      imemBusCtrl_commitValid <= 1'b0;
    end else begin
      if(when_VliwSimdSoc_l135) begin
        imemBusCtrl_bothFired <= 1'b1;
        imemBusCtrl_awDone <= 1'b0;
        imemBusCtrl_wDone <= 1'b0;
        imemBusCtrl_awReady <= 1'b0;
        imemBusCtrl_wReady <= 1'b0;
      end else begin
        if(imemBusCtrl_awFire) begin
          imemBusCtrl_awDone <= 1'b1;
          imemBusCtrl_awReady <= 1'b0;
        end else begin
          if(imemBusCtrl_wFire) begin
            imemBusCtrl_wDone <= 1'b1;
            imemBusCtrl_wReady <= 1'b0;
          end
        end
      end
      if(when_VliwSimdSoc_l149) begin
        imemBusCtrl_bothFired <= 1'b1;
        imemBusCtrl_awDone <= 1'b0;
        imemBusCtrl_wDone <= 1'b0;
        imemBusCtrl_awReady <= 1'b0;
        imemBusCtrl_wReady <= 1'b0;
      end
      if(when_VliwSimdSoc_l156) begin
        imemBusCtrl_bothFired <= 1'b1;
        imemBusCtrl_awDone <= 1'b0;
        imemBusCtrl_wDone <= 1'b0;
        imemBusCtrl_awReady <= 1'b0;
        imemBusCtrl_wReady <= 1'b0;
      end
      if(imemBusCtrl_bothFired) begin
        imemBusCtrl_accumulator[_zz_imemBusCtrl_accumulator_1] <= imemBusCtrl_wData[0];
        imemBusCtrl_accumulator[_zz_imemBusCtrl_accumulator_3] <= imemBusCtrl_wData[1];
        imemBusCtrl_accumulator[_zz_imemBusCtrl_accumulator_5] <= imemBusCtrl_wData[2];
        imemBusCtrl_accumulator[_zz_imemBusCtrl_accumulator_7] <= imemBusCtrl_wData[3];
        imemBusCtrl_accumulator[_zz_imemBusCtrl_accumulator_9] <= imemBusCtrl_wData[4];
        imemBusCtrl_accumulator[_zz_imemBusCtrl_accumulator_11] <= imemBusCtrl_wData[5];
        imemBusCtrl_accumulator[_zz_imemBusCtrl_accumulator_13] <= imemBusCtrl_wData[6];
        imemBusCtrl_accumulator[_zz_imemBusCtrl_accumulator_15] <= imemBusCtrl_wData[7];
        imemBusCtrl_accumulator[_zz_imemBusCtrl_accumulator_17] <= imemBusCtrl_wData[8];
        imemBusCtrl_accumulator[_zz_imemBusCtrl_accumulator_19] <= imemBusCtrl_wData[9];
        imemBusCtrl_accumulator[_zz_imemBusCtrl_accumulator_21] <= imemBusCtrl_wData[10];
        imemBusCtrl_accumulator[_zz_imemBusCtrl_accumulator_23] <= imemBusCtrl_wData[11];
        imemBusCtrl_accumulator[_zz_imemBusCtrl_accumulator_25] <= imemBusCtrl_wData[12];
        imemBusCtrl_accumulator[_zz_imemBusCtrl_accumulator_27] <= imemBusCtrl_wData[13];
        imemBusCtrl_accumulator[_zz_imemBusCtrl_accumulator_29] <= imemBusCtrl_wData[14];
        imemBusCtrl_accumulator[_zz_imemBusCtrl_accumulator_31] <= imemBusCtrl_wData[15];
        imemBusCtrl_accumulator[_zz_imemBusCtrl_accumulator_33] <= imemBusCtrl_wData[16];
        imemBusCtrl_accumulator[_zz_imemBusCtrl_accumulator_35] <= imemBusCtrl_wData[17];
        imemBusCtrl_accumulator[_zz_imemBusCtrl_accumulator_37] <= imemBusCtrl_wData[18];
        imemBusCtrl_accumulator[_zz_imemBusCtrl_accumulator_39] <= imemBusCtrl_wData[19];
        imemBusCtrl_accumulator[_zz_imemBusCtrl_accumulator_41] <= imemBusCtrl_wData[20];
        imemBusCtrl_accumulator[_zz_imemBusCtrl_accumulator_43] <= imemBusCtrl_wData[21];
        imemBusCtrl_accumulator[_zz_imemBusCtrl_accumulator_45] <= imemBusCtrl_wData[22];
        imemBusCtrl_accumulator[_zz_imemBusCtrl_accumulator_47] <= imemBusCtrl_wData[23];
        imemBusCtrl_accumulator[_zz_imemBusCtrl_accumulator_49] <= imemBusCtrl_wData[24];
        imemBusCtrl_accumulator[_zz_imemBusCtrl_accumulator_51] <= imemBusCtrl_wData[25];
        imemBusCtrl_accumulator[_zz_imemBusCtrl_accumulator_53] <= imemBusCtrl_wData[26];
        imemBusCtrl_accumulator[_zz_imemBusCtrl_accumulator_55] <= imemBusCtrl_wData[27];
        imemBusCtrl_accumulator[_zz_imemBusCtrl_accumulator_57] <= imemBusCtrl_wData[28];
        imemBusCtrl_accumulator[_zz_imemBusCtrl_accumulator_59] <= imemBusCtrl_wData[29];
        imemBusCtrl_accumulator[_zz_imemBusCtrl_accumulator_61] <= imemBusCtrl_wData[30];
        imemBusCtrl_accumulator[_zz_imemBusCtrl_accumulator_63] <= imemBusCtrl_wData[31];
      end
      imemBusCtrl_commitValid <= (imemBusCtrl_bothFired && imemBusCtrl_isLastWord);
      if(imemBusCtrl_bothFired) begin
        imemBusCtrl_bValid <= 1'b1;
      end
      if(when_VliwSimdSoc_l228) begin
        imemBusCtrl_bValid <= 1'b0;
        imemBusCtrl_awReady <= 1'b1;
        imemBusCtrl_wReady <= 1'b1;
        imemBusCtrl_bothFired <= 1'b0;
      end
    end
  end

  always @(posedge clk) begin
    if(imemBusCtrl_awFire) begin
      imemBusCtrl_awAddr <= io_imemAxi_aw_payload_addr;
    end
    if(imemBusCtrl_wFire) begin
      imemBusCtrl_wData <= io_imemAxi_w_payload_data;
    end
    imemBusCtrl_commitAddr <= imemBusCtrl_instrAddr;
    imemBusCtrl_commitCore <= imemBusCtrl_coreSelect;
    if(when_VliwSimdSoc_l204) begin
      imemBusCtrl_commitData <= imemBusCtrl_accumulator;
      imemBusCtrl_commitData[_zz_imemBusCtrl_commitData_1] <= imemBusCtrl_wData[0];
      imemBusCtrl_commitData[_zz_imemBusCtrl_commitData_3] <= imemBusCtrl_wData[1];
      imemBusCtrl_commitData[_zz_imemBusCtrl_commitData_5] <= imemBusCtrl_wData[2];
      imemBusCtrl_commitData[_zz_imemBusCtrl_commitData_7] <= imemBusCtrl_wData[3];
      imemBusCtrl_commitData[_zz_imemBusCtrl_commitData_9] <= imemBusCtrl_wData[4];
      imemBusCtrl_commitData[_zz_imemBusCtrl_commitData_11] <= imemBusCtrl_wData[5];
      imemBusCtrl_commitData[_zz_imemBusCtrl_commitData_13] <= imemBusCtrl_wData[6];
      imemBusCtrl_commitData[_zz_imemBusCtrl_commitData_15] <= imemBusCtrl_wData[7];
      imemBusCtrl_commitData[_zz_imemBusCtrl_commitData_17] <= imemBusCtrl_wData[8];
      imemBusCtrl_commitData[_zz_imemBusCtrl_commitData_19] <= imemBusCtrl_wData[9];
      imemBusCtrl_commitData[_zz_imemBusCtrl_commitData_21] <= imemBusCtrl_wData[10];
      imemBusCtrl_commitData[_zz_imemBusCtrl_commitData_23] <= imemBusCtrl_wData[11];
      imemBusCtrl_commitData[_zz_imemBusCtrl_commitData_25] <= imemBusCtrl_wData[12];
      imemBusCtrl_commitData[_zz_imemBusCtrl_commitData_27] <= imemBusCtrl_wData[13];
      imemBusCtrl_commitData[_zz_imemBusCtrl_commitData_29] <= imemBusCtrl_wData[14];
      imemBusCtrl_commitData[_zz_imemBusCtrl_commitData_31] <= imemBusCtrl_wData[15];
      imemBusCtrl_commitData[_zz_imemBusCtrl_commitData_33] <= imemBusCtrl_wData[16];
      imemBusCtrl_commitData[_zz_imemBusCtrl_commitData_35] <= imemBusCtrl_wData[17];
      imemBusCtrl_commitData[_zz_imemBusCtrl_commitData_37] <= imemBusCtrl_wData[18];
      imemBusCtrl_commitData[_zz_imemBusCtrl_commitData_39] <= imemBusCtrl_wData[19];
      imemBusCtrl_commitData[_zz_imemBusCtrl_commitData_41] <= imemBusCtrl_wData[20];
      imemBusCtrl_commitData[_zz_imemBusCtrl_commitData_43] <= imemBusCtrl_wData[21];
      imemBusCtrl_commitData[_zz_imemBusCtrl_commitData_45] <= imemBusCtrl_wData[22];
      imemBusCtrl_commitData[_zz_imemBusCtrl_commitData_47] <= imemBusCtrl_wData[23];
      imemBusCtrl_commitData[_zz_imemBusCtrl_commitData_49] <= imemBusCtrl_wData[24];
      imemBusCtrl_commitData[_zz_imemBusCtrl_commitData_51] <= imemBusCtrl_wData[25];
      imemBusCtrl_commitData[_zz_imemBusCtrl_commitData_53] <= imemBusCtrl_wData[26];
      imemBusCtrl_commitData[_zz_imemBusCtrl_commitData_55] <= imemBusCtrl_wData[27];
      imemBusCtrl_commitData[_zz_imemBusCtrl_commitData_57] <= imemBusCtrl_wData[28];
      imemBusCtrl_commitData[_zz_imemBusCtrl_commitData_59] <= imemBusCtrl_wData[29];
      imemBusCtrl_commitData[_zz_imemBusCtrl_commitData_61] <= imemBusCtrl_wData[30];
      imemBusCtrl_commitData[_zz_imemBusCtrl_commitData_63] <= imemBusCtrl_wData[31];
    end
  end


endmodule

module HostInterface (
  input  wire          io_axiLite_aw_valid,
  output wire          io_axiLite_aw_ready,
  input  wire [31:0]   io_axiLite_aw_payload_addr,
  input  wire [2:0]    io_axiLite_aw_payload_prot,
  input  wire          io_axiLite_w_valid,
  output wire          io_axiLite_w_ready,
  input  wire [31:0]   io_axiLite_w_payload_data,
  input  wire [3:0]    io_axiLite_w_payload_strb,
  output wire          io_axiLite_b_valid,
  input  wire          io_axiLite_b_ready,
  output wire [1:0]    io_axiLite_b_payload_resp,
  input  wire          io_axiLite_ar_valid,
  output wire          io_axiLite_ar_ready,
  input  wire [31:0]   io_axiLite_ar_payload_addr,
  input  wire [2:0]    io_axiLite_ar_payload_prot,
  output wire          io_axiLite_r_valid,
  input  wire          io_axiLite_r_ready,
  output wire [31:0]   io_axiLite_r_payload_data,
  output wire [1:0]    io_axiLite_r_payload_resp,
  output wire          io_coreStart_0,
  output wire          io_coreReset_0,
  input  wire          io_coreHalted_0,
  input  wire          io_coreRunning_0,
  input  wire [9:0]    io_corePc_0,
  input  wire [31:0]   io_coreCycles_0,
  output wire          io_irq,
  input  wire          clk,
  input  wire          reset
);

  wire       [31:0]   _zz_busCtrl_readRsp_data;
  wire                busCtrl_readErrorFlag;
  wire                busCtrl_writeErrorFlag;
  wire                busCtrl_readHaltRequest;
  wire                busCtrl_writeHaltRequest;
  wire                busCtrl_writeJoinEvent_valid;
  wire                busCtrl_writeJoinEvent_ready;
  wire                busCtrl_writeOccur;
  reg        [1:0]    busCtrl_writeRsp_resp;
  wire                busCtrl_writeJoinEvent_translated_valid;
  wire                busCtrl_writeJoinEvent_translated_ready;
  wire       [1:0]    busCtrl_writeJoinEvent_translated_payload_resp;
  wire                _zz_busCtrl_writeJoinEvent_translated_ready;
  wire                _zz_busCtrl_writeJoinEvent_translated_ready_1;
  wire                _zz_io_axiLite_b_valid;
  reg                 _zz_io_axiLite_b_valid_1;
  reg        [1:0]    _zz_io_axiLite_b_payload_resp;
  wire                busCtrl_readDataStage_valid;
  wire                busCtrl_readDataStage_ready;
  wire       [31:0]   busCtrl_readDataStage_payload_addr;
  wire       [2:0]    busCtrl_readDataStage_payload_prot;
  reg                 io_axiLite_ar_rValid;
  wire                busCtrl_readDataStage_fire;
  reg        [31:0]   io_axiLite_ar_rData_addr;
  reg        [2:0]    io_axiLite_ar_rData_prot;
  reg        [31:0]   busCtrl_readRsp_data;
  reg        [1:0]    busCtrl_readRsp_resp;
  wire                _zz_io_axiLite_r_valid;
  wire       [31:0]   busCtrl_readAddressMasked;
  wire       [31:0]   busCtrl_writeAddressMasked;
  wire                busCtrl_readOccur;
  reg        [31:0]   ctrlReg;
  reg                 _zz_startPulse;
  wire                startPulse;
  reg                 _zz_resetPulse;
  wire                resetPulse;
  reg        [31:0]   statusReg;
  reg        [31:0]   globalCycleCounter;
  reg        [31:0]   slotConfigBits;
  reg                 anyStarted;
  function [31:0] zz_slotConfigBits(input dummy);
    begin
      zz_slotConfigBits = 32'h0;
      zz_slotConfigBits[3 : 0] = 4'b0001;
      zz_slotConfigBits[7 : 4] = 4'b0001;
      zz_slotConfigBits[11 : 8] = 4'b0001;
      zz_slotConfigBits[15 : 12] = 4'b0001;
    end
  endfunction
  wire [31:0] _zz_1;

  assign _zz_busCtrl_readRsp_data = {22'd0, io_corePc_0};
  assign busCtrl_readErrorFlag = 1'b0;
  assign busCtrl_writeErrorFlag = 1'b0;
  assign busCtrl_readHaltRequest = 1'b0;
  assign busCtrl_writeHaltRequest = 1'b0;
  assign busCtrl_writeOccur = (busCtrl_writeJoinEvent_valid && busCtrl_writeJoinEvent_ready);
  assign busCtrl_writeJoinEvent_valid = (io_axiLite_aw_valid && io_axiLite_w_valid);
  assign io_axiLite_aw_ready = busCtrl_writeOccur;
  assign io_axiLite_w_ready = busCtrl_writeOccur;
  assign busCtrl_writeJoinEvent_translated_valid = busCtrl_writeJoinEvent_valid;
  assign busCtrl_writeJoinEvent_ready = busCtrl_writeJoinEvent_translated_ready;
  assign busCtrl_writeJoinEvent_translated_payload_resp = busCtrl_writeRsp_resp;
  assign _zz_busCtrl_writeJoinEvent_translated_ready = (! busCtrl_writeHaltRequest);
  assign busCtrl_writeJoinEvent_translated_ready = (_zz_busCtrl_writeJoinEvent_translated_ready_1 && _zz_busCtrl_writeJoinEvent_translated_ready);
  assign _zz_busCtrl_writeJoinEvent_translated_ready_1 = (! _zz_io_axiLite_b_valid_1);
  assign _zz_io_axiLite_b_valid = _zz_io_axiLite_b_valid_1;
  assign io_axiLite_b_valid = _zz_io_axiLite_b_valid;
  assign io_axiLite_b_payload_resp = _zz_io_axiLite_b_payload_resp;
  assign busCtrl_readDataStage_fire = (busCtrl_readDataStage_valid && busCtrl_readDataStage_ready);
  assign io_axiLite_ar_ready = (! io_axiLite_ar_rValid);
  assign busCtrl_readDataStage_valid = io_axiLite_ar_rValid;
  assign busCtrl_readDataStage_payload_addr = io_axiLite_ar_rData_addr;
  assign busCtrl_readDataStage_payload_prot = io_axiLite_ar_rData_prot;
  assign _zz_io_axiLite_r_valid = (! busCtrl_readHaltRequest);
  assign busCtrl_readDataStage_ready = (io_axiLite_r_ready && _zz_io_axiLite_r_valid);
  assign io_axiLite_r_valid = (busCtrl_readDataStage_valid && _zz_io_axiLite_r_valid);
  assign io_axiLite_r_payload_data = busCtrl_readRsp_data;
  assign io_axiLite_r_payload_resp = busCtrl_readRsp_resp;
  always @(*) begin
    if(busCtrl_writeErrorFlag) begin
      busCtrl_writeRsp_resp = 2'b10;
    end else begin
      busCtrl_writeRsp_resp = 2'b00;
    end
  end

  always @(*) begin
    if(busCtrl_readErrorFlag) begin
      busCtrl_readRsp_resp = 2'b10;
    end else begin
      busCtrl_readRsp_resp = 2'b00;
    end
  end

  always @(*) begin
    busCtrl_readRsp_data = 32'h0;
    case(busCtrl_readAddressMasked)
      32'h0 : begin
        busCtrl_readRsp_data[31 : 0] = ctrlReg;
      end
      32'h00000004 : begin
        busCtrl_readRsp_data[31 : 0] = statusReg;
      end
      32'h00000008 : begin
        busCtrl_readRsp_data[31 : 0] = globalCycleCounter;
      end
      32'h0000000c : begin
        busCtrl_readRsp_data[31 : 0] = 32'h00000001;
      end
      32'h00000010 : begin
        busCtrl_readRsp_data[31 : 0] = 32'h00000008;
      end
      32'h00000014 : begin
        busCtrl_readRsp_data[31 : 0] = 32'h00000600;
      end
      32'h00000018 : begin
        busCtrl_readRsp_data[31 : 0] = 32'h00000400;
      end
      32'h0000001c : begin
        busCtrl_readRsp_data[31 : 0] = 32'h00000100;
      end
      32'h00000020 : begin
        busCtrl_readRsp_data[31 : 0] = slotConfigBits;
      end
      32'h00000100 : begin
        busCtrl_readRsp_data[31 : 0] = _zz_busCtrl_readRsp_data;
      end
      32'h00000200 : begin
        busCtrl_readRsp_data[31 : 0] = io_coreCycles_0;
      end
      default : begin
      end
    endcase
  end

  assign busCtrl_readAddressMasked = (busCtrl_readDataStage_payload_addr & (~ 32'h00000003));
  assign busCtrl_writeAddressMasked = (io_axiLite_aw_payload_addr & (~ 32'h00000003));
  assign busCtrl_readOccur = (io_axiLite_r_valid && io_axiLite_r_ready);
  assign startPulse = (ctrlReg[0] && (! _zz_startPulse));
  assign resetPulse = (ctrlReg[1] && (! _zz_resetPulse));
  assign io_coreStart_0 = startPulse;
  assign io_coreReset_0 = resetPulse;
  always @(*) begin
    statusReg = 32'h0;
    statusReg[0] = io_coreRunning_0;
    statusReg[1] = io_coreHalted_0;
  end

  assign _zz_1 = zz_slotConfigBits(1'b0);
  always @(*) slotConfigBits = _zz_1;
  assign io_irq = (anyStarted && io_coreHalted_0);
  always @(posedge clk) begin
    if(reset) begin
      _zz_io_axiLite_b_valid_1 <= 1'b0;
      io_axiLite_ar_rValid <= 1'b0;
      ctrlReg <= 32'h0;
      _zz_startPulse <= 1'b0;
      _zz_resetPulse <= 1'b0;
      globalCycleCounter <= 32'h0;
      anyStarted <= 1'b0;
    end else begin
      if((busCtrl_writeJoinEvent_translated_valid && _zz_busCtrl_writeJoinEvent_translated_ready)) begin
        _zz_io_axiLite_b_valid_1 <= 1'b1;
      end
      if((_zz_io_axiLite_b_valid && io_axiLite_b_ready)) begin
        _zz_io_axiLite_b_valid_1 <= 1'b0;
      end
      if(io_axiLite_ar_valid) begin
        io_axiLite_ar_rValid <= 1'b1;
      end
      if(busCtrl_readDataStage_fire) begin
        io_axiLite_ar_rValid <= 1'b0;
      end
      _zz_startPulse <= ctrlReg[0];
      _zz_resetPulse <= ctrlReg[1];
      if(startPulse) begin
        ctrlReg[0] <= 1'b0;
      end
      if(resetPulse) begin
        ctrlReg[1] <= 1'b0;
      end
      if(io_coreRunning_0) begin
        globalCycleCounter <= (globalCycleCounter + 32'h00000001);
      end
      if(startPulse) begin
        anyStarted <= 1'b1;
      end
      if(resetPulse) begin
        anyStarted <= 1'b0;
      end
      case(busCtrl_writeAddressMasked)
        32'h0 : begin
          if(busCtrl_writeOccur) begin
            ctrlReg <= io_axiLite_w_payload_data[31 : 0];
          end
        end
        default : begin
        end
      endcase
    end
  end

  always @(posedge clk) begin
    if(_zz_busCtrl_writeJoinEvent_translated_ready_1) begin
      _zz_io_axiLite_b_payload_resp <= busCtrl_writeJoinEvent_translated_payload_resp;
    end
    if(io_axiLite_ar_ready) begin
      io_axiLite_ar_rData_addr <= io_axiLite_ar_payload_addr;
      io_axiLite_ar_rData_prot <= io_axiLite_ar_payload_prot;
    end
  end


endmodule

module MemorySubsystem (
  input  wire          io_corePorts_0_aw_valid,
  output wire          io_corePorts_0_aw_ready,
  input  wire [31:0]   io_corePorts_0_aw_payload_addr,
  input  wire [3:0]    io_corePorts_0_aw_payload_id,
  input  wire [7:0]    io_corePorts_0_aw_payload_len,
  input  wire [2:0]    io_corePorts_0_aw_payload_size,
  input  wire [1:0]    io_corePorts_0_aw_payload_burst,
  input  wire          io_corePorts_0_w_valid,
  output wire          io_corePorts_0_w_ready,
  input  wire [31:0]   io_corePorts_0_w_payload_data,
  input  wire [3:0]    io_corePorts_0_w_payload_strb,
  input  wire          io_corePorts_0_w_payload_last,
  output wire          io_corePorts_0_b_valid,
  input  wire          io_corePorts_0_b_ready,
  output wire [3:0]    io_corePorts_0_b_payload_id,
  output wire [1:0]    io_corePorts_0_b_payload_resp,
  input  wire          io_corePorts_0_ar_valid,
  output wire          io_corePorts_0_ar_ready,
  input  wire [31:0]   io_corePorts_0_ar_payload_addr,
  input  wire [3:0]    io_corePorts_0_ar_payload_id,
  input  wire [7:0]    io_corePorts_0_ar_payload_len,
  input  wire [2:0]    io_corePorts_0_ar_payload_size,
  input  wire [1:0]    io_corePorts_0_ar_payload_burst,
  output wire          io_corePorts_0_r_valid,
  input  wire          io_corePorts_0_r_ready,
  output wire [31:0]   io_corePorts_0_r_payload_data,
  output wire [3:0]    io_corePorts_0_r_payload_id,
  output wire [1:0]    io_corePorts_0_r_payload_resp,
  output wire          io_corePorts_0_r_payload_last,
  input  wire          io_hostPort_aw_valid,
  output wire          io_hostPort_aw_ready,
  input  wire [31:0]   io_hostPort_aw_payload_addr,
  input  wire [3:0]    io_hostPort_aw_payload_id,
  input  wire [7:0]    io_hostPort_aw_payload_len,
  input  wire [2:0]    io_hostPort_aw_payload_size,
  input  wire [1:0]    io_hostPort_aw_payload_burst,
  input  wire          io_hostPort_w_valid,
  output wire          io_hostPort_w_ready,
  input  wire [31:0]   io_hostPort_w_payload_data,
  input  wire [3:0]    io_hostPort_w_payload_strb,
  input  wire          io_hostPort_w_payload_last,
  output wire          io_hostPort_b_valid,
  input  wire          io_hostPort_b_ready,
  output wire [3:0]    io_hostPort_b_payload_id,
  output wire [1:0]    io_hostPort_b_payload_resp,
  input  wire          io_hostPort_ar_valid,
  output wire          io_hostPort_ar_ready,
  input  wire [31:0]   io_hostPort_ar_payload_addr,
  input  wire [3:0]    io_hostPort_ar_payload_id,
  input  wire [7:0]    io_hostPort_ar_payload_len,
  input  wire [2:0]    io_hostPort_ar_payload_size,
  input  wire [1:0]    io_hostPort_ar_payload_burst,
  output wire          io_hostPort_r_valid,
  input  wire          io_hostPort_r_ready,
  output wire [31:0]   io_hostPort_r_payload_data,
  output wire [3:0]    io_hostPort_r_payload_id,
  output wire [1:0]    io_hostPort_r_payload_resp,
  output wire          io_hostPort_r_payload_last,
  input  wire          clk,
  input  wire          reset
);

  wire       [3:0]    io_corePorts_0_readOnly_decoder_io_outputs_0_r_payload_id;
  wire       [3:0]    io_corePorts_0_writeOnly_decoder_io_outputs_0_b_payload_id;
  wire       [3:0]    io_hostPort_readOnly_decoder_io_outputs_0_r_payload_id;
  wire       [3:0]    io_hostPort_writeOnly_decoder_io_outputs_0_b_payload_id;
  wire       [15:0]   ram_io_axi_arbiter_io_readInputs_0_ar_payload_addr;
  wire       [4:0]    ram_io_axi_arbiter_io_readInputs_0_ar_payload_id;
  wire       [15:0]   ram_io_axi_arbiter_io_readInputs_1_ar_payload_addr;
  wire       [4:0]    ram_io_axi_arbiter_io_readInputs_1_ar_payload_id;
  wire       [15:0]   ram_io_axi_arbiter_io_writeInputs_0_aw_payload_addr;
  wire       [4:0]    ram_io_axi_arbiter_io_writeInputs_0_aw_payload_id;
  wire       [15:0]   ram_io_axi_arbiter_io_writeInputs_1_aw_payload_addr;
  wire       [4:0]    ram_io_axi_arbiter_io_writeInputs_1_aw_payload_id;
  wire                ram_io_axi_arw_ready;
  wire                ram_io_axi_w_ready;
  wire                ram_io_axi_b_valid;
  wire       [5:0]    ram_io_axi_b_payload_id;
  wire       [1:0]    ram_io_axi_b_payload_resp;
  wire                ram_io_axi_r_valid;
  wire       [31:0]   ram_io_axi_r_payload_data;
  wire       [5:0]    ram_io_axi_r_payload_id;
  wire       [1:0]    ram_io_axi_r_payload_resp;
  wire                ram_io_axi_r_payload_last;
  wire                io_corePorts_0_readOnly_decoder_io_input_ar_ready;
  wire                io_corePorts_0_readOnly_decoder_io_input_r_valid;
  wire       [31:0]   io_corePorts_0_readOnly_decoder_io_input_r_payload_data;
  wire       [3:0]    io_corePorts_0_readOnly_decoder_io_input_r_payload_id;
  wire       [1:0]    io_corePorts_0_readOnly_decoder_io_input_r_payload_resp;
  wire                io_corePorts_0_readOnly_decoder_io_input_r_payload_last;
  wire                io_corePorts_0_readOnly_decoder_io_outputs_0_ar_valid;
  wire       [31:0]   io_corePorts_0_readOnly_decoder_io_outputs_0_ar_payload_addr;
  wire       [3:0]    io_corePorts_0_readOnly_decoder_io_outputs_0_ar_payload_id;
  wire       [7:0]    io_corePorts_0_readOnly_decoder_io_outputs_0_ar_payload_len;
  wire       [2:0]    io_corePorts_0_readOnly_decoder_io_outputs_0_ar_payload_size;
  wire       [1:0]    io_corePorts_0_readOnly_decoder_io_outputs_0_ar_payload_burst;
  wire                io_corePorts_0_readOnly_decoder_io_outputs_0_r_ready;
  wire                io_corePorts_0_writeOnly_decoder_io_input_aw_ready;
  wire                io_corePorts_0_writeOnly_decoder_io_input_w_ready;
  wire                io_corePorts_0_writeOnly_decoder_io_input_b_valid;
  wire       [3:0]    io_corePorts_0_writeOnly_decoder_io_input_b_payload_id;
  wire       [1:0]    io_corePorts_0_writeOnly_decoder_io_input_b_payload_resp;
  wire                io_corePorts_0_writeOnly_decoder_io_outputs_0_aw_valid;
  wire       [31:0]   io_corePorts_0_writeOnly_decoder_io_outputs_0_aw_payload_addr;
  wire       [3:0]    io_corePorts_0_writeOnly_decoder_io_outputs_0_aw_payload_id;
  wire       [7:0]    io_corePorts_0_writeOnly_decoder_io_outputs_0_aw_payload_len;
  wire       [2:0]    io_corePorts_0_writeOnly_decoder_io_outputs_0_aw_payload_size;
  wire       [1:0]    io_corePorts_0_writeOnly_decoder_io_outputs_0_aw_payload_burst;
  wire                io_corePorts_0_writeOnly_decoder_io_outputs_0_w_valid;
  wire       [31:0]   io_corePorts_0_writeOnly_decoder_io_outputs_0_w_payload_data;
  wire       [3:0]    io_corePorts_0_writeOnly_decoder_io_outputs_0_w_payload_strb;
  wire                io_corePorts_0_writeOnly_decoder_io_outputs_0_w_payload_last;
  wire                io_corePorts_0_writeOnly_decoder_io_outputs_0_b_ready;
  wire                io_hostPort_readOnly_decoder_io_input_ar_ready;
  wire                io_hostPort_readOnly_decoder_io_input_r_valid;
  wire       [31:0]   io_hostPort_readOnly_decoder_io_input_r_payload_data;
  wire       [3:0]    io_hostPort_readOnly_decoder_io_input_r_payload_id;
  wire       [1:0]    io_hostPort_readOnly_decoder_io_input_r_payload_resp;
  wire                io_hostPort_readOnly_decoder_io_input_r_payload_last;
  wire                io_hostPort_readOnly_decoder_io_outputs_0_ar_valid;
  wire       [31:0]   io_hostPort_readOnly_decoder_io_outputs_0_ar_payload_addr;
  wire       [3:0]    io_hostPort_readOnly_decoder_io_outputs_0_ar_payload_id;
  wire       [7:0]    io_hostPort_readOnly_decoder_io_outputs_0_ar_payload_len;
  wire       [2:0]    io_hostPort_readOnly_decoder_io_outputs_0_ar_payload_size;
  wire       [1:0]    io_hostPort_readOnly_decoder_io_outputs_0_ar_payload_burst;
  wire                io_hostPort_readOnly_decoder_io_outputs_0_r_ready;
  wire                io_hostPort_writeOnly_decoder_io_input_aw_ready;
  wire                io_hostPort_writeOnly_decoder_io_input_w_ready;
  wire                io_hostPort_writeOnly_decoder_io_input_b_valid;
  wire       [3:0]    io_hostPort_writeOnly_decoder_io_input_b_payload_id;
  wire       [1:0]    io_hostPort_writeOnly_decoder_io_input_b_payload_resp;
  wire                io_hostPort_writeOnly_decoder_io_outputs_0_aw_valid;
  wire       [31:0]   io_hostPort_writeOnly_decoder_io_outputs_0_aw_payload_addr;
  wire       [3:0]    io_hostPort_writeOnly_decoder_io_outputs_0_aw_payload_id;
  wire       [7:0]    io_hostPort_writeOnly_decoder_io_outputs_0_aw_payload_len;
  wire       [2:0]    io_hostPort_writeOnly_decoder_io_outputs_0_aw_payload_size;
  wire       [1:0]    io_hostPort_writeOnly_decoder_io_outputs_0_aw_payload_burst;
  wire                io_hostPort_writeOnly_decoder_io_outputs_0_w_valid;
  wire       [31:0]   io_hostPort_writeOnly_decoder_io_outputs_0_w_payload_data;
  wire       [3:0]    io_hostPort_writeOnly_decoder_io_outputs_0_w_payload_strb;
  wire                io_hostPort_writeOnly_decoder_io_outputs_0_w_payload_last;
  wire                io_hostPort_writeOnly_decoder_io_outputs_0_b_ready;
  wire                ram_io_axi_arbiter_io_readInputs_0_ar_ready;
  wire                ram_io_axi_arbiter_io_readInputs_0_r_valid;
  wire       [31:0]   ram_io_axi_arbiter_io_readInputs_0_r_payload_data;
  wire       [4:0]    ram_io_axi_arbiter_io_readInputs_0_r_payload_id;
  wire       [1:0]    ram_io_axi_arbiter_io_readInputs_0_r_payload_resp;
  wire                ram_io_axi_arbiter_io_readInputs_0_r_payload_last;
  wire                ram_io_axi_arbiter_io_readInputs_1_ar_ready;
  wire                ram_io_axi_arbiter_io_readInputs_1_r_valid;
  wire       [31:0]   ram_io_axi_arbiter_io_readInputs_1_r_payload_data;
  wire       [4:0]    ram_io_axi_arbiter_io_readInputs_1_r_payload_id;
  wire       [1:0]    ram_io_axi_arbiter_io_readInputs_1_r_payload_resp;
  wire                ram_io_axi_arbiter_io_readInputs_1_r_payload_last;
  wire                ram_io_axi_arbiter_io_writeInputs_0_aw_ready;
  wire                ram_io_axi_arbiter_io_writeInputs_0_w_ready;
  wire                ram_io_axi_arbiter_io_writeInputs_0_b_valid;
  wire       [4:0]    ram_io_axi_arbiter_io_writeInputs_0_b_payload_id;
  wire       [1:0]    ram_io_axi_arbiter_io_writeInputs_0_b_payload_resp;
  wire                ram_io_axi_arbiter_io_writeInputs_1_aw_ready;
  wire                ram_io_axi_arbiter_io_writeInputs_1_w_ready;
  wire                ram_io_axi_arbiter_io_writeInputs_1_b_valid;
  wire       [4:0]    ram_io_axi_arbiter_io_writeInputs_1_b_payload_id;
  wire       [1:0]    ram_io_axi_arbiter_io_writeInputs_1_b_payload_resp;
  wire                ram_io_axi_arbiter_io_output_arw_valid;
  wire       [15:0]   ram_io_axi_arbiter_io_output_arw_payload_addr;
  wire       [5:0]    ram_io_axi_arbiter_io_output_arw_payload_id;
  wire       [7:0]    ram_io_axi_arbiter_io_output_arw_payload_len;
  wire       [2:0]    ram_io_axi_arbiter_io_output_arw_payload_size;
  wire       [1:0]    ram_io_axi_arbiter_io_output_arw_payload_burst;
  wire                ram_io_axi_arbiter_io_output_arw_payload_write;
  wire                ram_io_axi_arbiter_io_output_w_valid;
  wire       [31:0]   ram_io_axi_arbiter_io_output_w_payload_data;
  wire       [3:0]    ram_io_axi_arbiter_io_output_w_payload_strb;
  wire                ram_io_axi_arbiter_io_output_w_payload_last;
  wire                ram_io_axi_arbiter_io_output_b_ready;
  wire                ram_io_axi_arbiter_io_output_r_ready;
  wire                io_corePorts_0_readOnly_ar_valid;
  wire                io_corePorts_0_readOnly_ar_ready;
  wire       [31:0]   io_corePorts_0_readOnly_ar_payload_addr;
  wire       [3:0]    io_corePorts_0_readOnly_ar_payload_id;
  wire       [7:0]    io_corePorts_0_readOnly_ar_payload_len;
  wire       [2:0]    io_corePorts_0_readOnly_ar_payload_size;
  wire       [1:0]    io_corePorts_0_readOnly_ar_payload_burst;
  wire                io_corePorts_0_readOnly_r_valid;
  wire                io_corePorts_0_readOnly_r_ready;
  wire       [31:0]   io_corePorts_0_readOnly_r_payload_data;
  wire       [3:0]    io_corePorts_0_readOnly_r_payload_id;
  wire       [1:0]    io_corePorts_0_readOnly_r_payload_resp;
  wire                io_corePorts_0_readOnly_r_payload_last;
  wire                io_corePorts_0_writeOnly_aw_valid;
  wire                io_corePorts_0_writeOnly_aw_ready;
  wire       [31:0]   io_corePorts_0_writeOnly_aw_payload_addr;
  wire       [3:0]    io_corePorts_0_writeOnly_aw_payload_id;
  wire       [7:0]    io_corePorts_0_writeOnly_aw_payload_len;
  wire       [2:0]    io_corePorts_0_writeOnly_aw_payload_size;
  wire       [1:0]    io_corePorts_0_writeOnly_aw_payload_burst;
  wire                io_corePorts_0_writeOnly_w_valid;
  wire                io_corePorts_0_writeOnly_w_ready;
  wire       [31:0]   io_corePorts_0_writeOnly_w_payload_data;
  wire       [3:0]    io_corePorts_0_writeOnly_w_payload_strb;
  wire                io_corePorts_0_writeOnly_w_payload_last;
  wire                io_corePorts_0_writeOnly_b_valid;
  wire                io_corePorts_0_writeOnly_b_ready;
  wire       [3:0]    io_corePorts_0_writeOnly_b_payload_id;
  wire       [1:0]    io_corePorts_0_writeOnly_b_payload_resp;
  wire                io_hostPort_readOnly_ar_valid;
  wire                io_hostPort_readOnly_ar_ready;
  wire       [31:0]   io_hostPort_readOnly_ar_payload_addr;
  wire       [3:0]    io_hostPort_readOnly_ar_payload_id;
  wire       [7:0]    io_hostPort_readOnly_ar_payload_len;
  wire       [2:0]    io_hostPort_readOnly_ar_payload_size;
  wire       [1:0]    io_hostPort_readOnly_ar_payload_burst;
  wire                io_hostPort_readOnly_r_valid;
  wire                io_hostPort_readOnly_r_ready;
  wire       [31:0]   io_hostPort_readOnly_r_payload_data;
  wire       [3:0]    io_hostPort_readOnly_r_payload_id;
  wire       [1:0]    io_hostPort_readOnly_r_payload_resp;
  wire                io_hostPort_readOnly_r_payload_last;
  wire                io_hostPort_writeOnly_aw_valid;
  wire                io_hostPort_writeOnly_aw_ready;
  wire       [31:0]   io_hostPort_writeOnly_aw_payload_addr;
  wire       [3:0]    io_hostPort_writeOnly_aw_payload_id;
  wire       [7:0]    io_hostPort_writeOnly_aw_payload_len;
  wire       [2:0]    io_hostPort_writeOnly_aw_payload_size;
  wire       [1:0]    io_hostPort_writeOnly_aw_payload_burst;
  wire                io_hostPort_writeOnly_w_valid;
  wire                io_hostPort_writeOnly_w_ready;
  wire       [31:0]   io_hostPort_writeOnly_w_payload_data;
  wire       [3:0]    io_hostPort_writeOnly_w_payload_strb;
  wire                io_hostPort_writeOnly_w_payload_last;
  wire                io_hostPort_writeOnly_b_valid;
  wire                io_hostPort_writeOnly_b_ready;
  wire       [3:0]    io_hostPort_writeOnly_b_payload_id;
  wire       [1:0]    io_hostPort_writeOnly_b_payload_resp;
  wire                memSub_io_corePorts_0_readOnly_decoder_io_outputs_0_ar_validPipe_valid;
  wire                memSub_io_corePorts_0_readOnly_decoder_io_outputs_0_ar_validPipe_ready;
  wire       [31:0]   memSub_io_corePorts_0_readOnly_decoder_io_outputs_0_ar_validPipe_payload_addr;
  wire       [3:0]    memSub_io_corePorts_0_readOnly_decoder_io_outputs_0_ar_validPipe_payload_id;
  wire       [7:0]    memSub_io_corePorts_0_readOnly_decoder_io_outputs_0_ar_validPipe_payload_len;
  wire       [2:0]    memSub_io_corePorts_0_readOnly_decoder_io_outputs_0_ar_validPipe_payload_size;
  wire       [1:0]    memSub_io_corePorts_0_readOnly_decoder_io_outputs_0_ar_validPipe_payload_burst;
  reg                 memSub_io_corePorts_0_readOnly_decoder_io_outputs_0_ar_rValid;
  wire                memSub_io_corePorts_0_readOnly_decoder_io_outputs_0_ar_validPipe_fire;
  wire                memSub_io_corePorts_0_writeOnly_decoder_io_outputs_0_aw_validPipe_valid;
  wire                memSub_io_corePorts_0_writeOnly_decoder_io_outputs_0_aw_validPipe_ready;
  wire       [31:0]   memSub_io_corePorts_0_writeOnly_decoder_io_outputs_0_aw_validPipe_payload_addr;
  wire       [3:0]    memSub_io_corePorts_0_writeOnly_decoder_io_outputs_0_aw_validPipe_payload_id;
  wire       [7:0]    memSub_io_corePorts_0_writeOnly_decoder_io_outputs_0_aw_validPipe_payload_len;
  wire       [2:0]    memSub_io_corePorts_0_writeOnly_decoder_io_outputs_0_aw_validPipe_payload_size;
  wire       [1:0]    memSub_io_corePorts_0_writeOnly_decoder_io_outputs_0_aw_validPipe_payload_burst;
  reg                 memSub_io_corePorts_0_writeOnly_decoder_io_outputs_0_aw_rValid;
  wire                memSub_io_corePorts_0_writeOnly_decoder_io_outputs_0_aw_validPipe_fire;
  wire                memSub_io_hostPort_readOnly_decoder_io_outputs_0_ar_validPipe_valid;
  wire                memSub_io_hostPort_readOnly_decoder_io_outputs_0_ar_validPipe_ready;
  wire       [31:0]   memSub_io_hostPort_readOnly_decoder_io_outputs_0_ar_validPipe_payload_addr;
  wire       [3:0]    memSub_io_hostPort_readOnly_decoder_io_outputs_0_ar_validPipe_payload_id;
  wire       [7:0]    memSub_io_hostPort_readOnly_decoder_io_outputs_0_ar_validPipe_payload_len;
  wire       [2:0]    memSub_io_hostPort_readOnly_decoder_io_outputs_0_ar_validPipe_payload_size;
  wire       [1:0]    memSub_io_hostPort_readOnly_decoder_io_outputs_0_ar_validPipe_payload_burst;
  reg                 memSub_io_hostPort_readOnly_decoder_io_outputs_0_ar_rValid;
  wire                memSub_io_hostPort_readOnly_decoder_io_outputs_0_ar_validPipe_fire;
  wire                memSub_io_hostPort_writeOnly_decoder_io_outputs_0_aw_validPipe_valid;
  wire                memSub_io_hostPort_writeOnly_decoder_io_outputs_0_aw_validPipe_ready;
  wire       [31:0]   memSub_io_hostPort_writeOnly_decoder_io_outputs_0_aw_validPipe_payload_addr;
  wire       [3:0]    memSub_io_hostPort_writeOnly_decoder_io_outputs_0_aw_validPipe_payload_id;
  wire       [7:0]    memSub_io_hostPort_writeOnly_decoder_io_outputs_0_aw_validPipe_payload_len;
  wire       [2:0]    memSub_io_hostPort_writeOnly_decoder_io_outputs_0_aw_validPipe_payload_size;
  wire       [1:0]    memSub_io_hostPort_writeOnly_decoder_io_outputs_0_aw_validPipe_payload_burst;
  reg                 memSub_io_hostPort_writeOnly_decoder_io_outputs_0_aw_rValid;
  wire                memSub_io_hostPort_writeOnly_decoder_io_outputs_0_aw_validPipe_fire;

  Axi4SharedOnChipRam ram (
    .io_axi_arw_valid         (ram_io_axi_arbiter_io_output_arw_valid             ), //i
    .io_axi_arw_ready         (ram_io_axi_arw_ready                               ), //o
    .io_axi_arw_payload_addr  (ram_io_axi_arbiter_io_output_arw_payload_addr[15:0]), //i
    .io_axi_arw_payload_id    (ram_io_axi_arbiter_io_output_arw_payload_id[5:0]   ), //i
    .io_axi_arw_payload_len   (ram_io_axi_arbiter_io_output_arw_payload_len[7:0]  ), //i
    .io_axi_arw_payload_size  (ram_io_axi_arbiter_io_output_arw_payload_size[2:0] ), //i
    .io_axi_arw_payload_burst (ram_io_axi_arbiter_io_output_arw_payload_burst[1:0]), //i
    .io_axi_arw_payload_write (ram_io_axi_arbiter_io_output_arw_payload_write     ), //i
    .io_axi_w_valid           (ram_io_axi_arbiter_io_output_w_valid               ), //i
    .io_axi_w_ready           (ram_io_axi_w_ready                                 ), //o
    .io_axi_w_payload_data    (ram_io_axi_arbiter_io_output_w_payload_data[31:0]  ), //i
    .io_axi_w_payload_strb    (ram_io_axi_arbiter_io_output_w_payload_strb[3:0]   ), //i
    .io_axi_w_payload_last    (ram_io_axi_arbiter_io_output_w_payload_last        ), //i
    .io_axi_b_valid           (ram_io_axi_b_valid                                 ), //o
    .io_axi_b_ready           (ram_io_axi_arbiter_io_output_b_ready               ), //i
    .io_axi_b_payload_id      (ram_io_axi_b_payload_id[5:0]                       ), //o
    .io_axi_b_payload_resp    (ram_io_axi_b_payload_resp[1:0]                     ), //o
    .io_axi_r_valid           (ram_io_axi_r_valid                                 ), //o
    .io_axi_r_ready           (ram_io_axi_arbiter_io_output_r_ready               ), //i
    .io_axi_r_payload_data    (ram_io_axi_r_payload_data[31:0]                    ), //o
    .io_axi_r_payload_id      (ram_io_axi_r_payload_id[5:0]                       ), //o
    .io_axi_r_payload_resp    (ram_io_axi_r_payload_resp[1:0]                     ), //o
    .io_axi_r_payload_last    (ram_io_axi_r_payload_last                          ), //o
    .clk                      (clk                                                ), //i
    .reset                    (reset                                              )  //i
  );
  Axi4ReadOnlyDecoder io_corePorts_0_readOnly_decoder (
    .io_input_ar_valid             (io_corePorts_0_readOnly_ar_valid                                     ), //i
    .io_input_ar_ready             (io_corePorts_0_readOnly_decoder_io_input_ar_ready                    ), //o
    .io_input_ar_payload_addr      (io_corePorts_0_readOnly_ar_payload_addr[31:0]                        ), //i
    .io_input_ar_payload_id        (io_corePorts_0_readOnly_ar_payload_id[3:0]                           ), //i
    .io_input_ar_payload_len       (io_corePorts_0_readOnly_ar_payload_len[7:0]                          ), //i
    .io_input_ar_payload_size      (io_corePorts_0_readOnly_ar_payload_size[2:0]                         ), //i
    .io_input_ar_payload_burst     (io_corePorts_0_readOnly_ar_payload_burst[1:0]                        ), //i
    .io_input_r_valid              (io_corePorts_0_readOnly_decoder_io_input_r_valid                     ), //o
    .io_input_r_ready              (io_corePorts_0_readOnly_r_ready                                      ), //i
    .io_input_r_payload_data       (io_corePorts_0_readOnly_decoder_io_input_r_payload_data[31:0]        ), //o
    .io_input_r_payload_id         (io_corePorts_0_readOnly_decoder_io_input_r_payload_id[3:0]           ), //o
    .io_input_r_payload_resp       (io_corePorts_0_readOnly_decoder_io_input_r_payload_resp[1:0]         ), //o
    .io_input_r_payload_last       (io_corePorts_0_readOnly_decoder_io_input_r_payload_last              ), //o
    .io_outputs_0_ar_valid         (io_corePorts_0_readOnly_decoder_io_outputs_0_ar_valid                ), //o
    .io_outputs_0_ar_ready         (memSub_io_corePorts_0_readOnly_decoder_io_outputs_0_ar_validPipe_fire), //i
    .io_outputs_0_ar_payload_addr  (io_corePorts_0_readOnly_decoder_io_outputs_0_ar_payload_addr[31:0]   ), //o
    .io_outputs_0_ar_payload_id    (io_corePorts_0_readOnly_decoder_io_outputs_0_ar_payload_id[3:0]      ), //o
    .io_outputs_0_ar_payload_len   (io_corePorts_0_readOnly_decoder_io_outputs_0_ar_payload_len[7:0]     ), //o
    .io_outputs_0_ar_payload_size  (io_corePorts_0_readOnly_decoder_io_outputs_0_ar_payload_size[2:0]    ), //o
    .io_outputs_0_ar_payload_burst (io_corePorts_0_readOnly_decoder_io_outputs_0_ar_payload_burst[1:0]   ), //o
    .io_outputs_0_r_valid          (ram_io_axi_arbiter_io_readInputs_0_r_valid                           ), //i
    .io_outputs_0_r_ready          (io_corePorts_0_readOnly_decoder_io_outputs_0_r_ready                 ), //o
    .io_outputs_0_r_payload_data   (ram_io_axi_arbiter_io_readInputs_0_r_payload_data[31:0]              ), //i
    .io_outputs_0_r_payload_id     (io_corePorts_0_readOnly_decoder_io_outputs_0_r_payload_id[3:0]       ), //i
    .io_outputs_0_r_payload_resp   (ram_io_axi_arbiter_io_readInputs_0_r_payload_resp[1:0]               ), //i
    .io_outputs_0_r_payload_last   (ram_io_axi_arbiter_io_readInputs_0_r_payload_last                    ), //i
    .clk                           (clk                                                                  ), //i
    .reset                         (reset                                                                )  //i
  );
  Axi4WriteOnlyDecoder io_corePorts_0_writeOnly_decoder (
    .io_input_aw_valid             (io_corePorts_0_writeOnly_aw_valid                                     ), //i
    .io_input_aw_ready             (io_corePorts_0_writeOnly_decoder_io_input_aw_ready                    ), //o
    .io_input_aw_payload_addr      (io_corePorts_0_writeOnly_aw_payload_addr[31:0]                        ), //i
    .io_input_aw_payload_id        (io_corePorts_0_writeOnly_aw_payload_id[3:0]                           ), //i
    .io_input_aw_payload_len       (io_corePorts_0_writeOnly_aw_payload_len[7:0]                          ), //i
    .io_input_aw_payload_size      (io_corePorts_0_writeOnly_aw_payload_size[2:0]                         ), //i
    .io_input_aw_payload_burst     (io_corePorts_0_writeOnly_aw_payload_burst[1:0]                        ), //i
    .io_input_w_valid              (io_corePorts_0_writeOnly_w_valid                                      ), //i
    .io_input_w_ready              (io_corePorts_0_writeOnly_decoder_io_input_w_ready                     ), //o
    .io_input_w_payload_data       (io_corePorts_0_writeOnly_w_payload_data[31:0]                         ), //i
    .io_input_w_payload_strb       (io_corePorts_0_writeOnly_w_payload_strb[3:0]                          ), //i
    .io_input_w_payload_last       (io_corePorts_0_writeOnly_w_payload_last                               ), //i
    .io_input_b_valid              (io_corePorts_0_writeOnly_decoder_io_input_b_valid                     ), //o
    .io_input_b_ready              (io_corePorts_0_writeOnly_b_ready                                      ), //i
    .io_input_b_payload_id         (io_corePorts_0_writeOnly_decoder_io_input_b_payload_id[3:0]           ), //o
    .io_input_b_payload_resp       (io_corePorts_0_writeOnly_decoder_io_input_b_payload_resp[1:0]         ), //o
    .io_outputs_0_aw_valid         (io_corePorts_0_writeOnly_decoder_io_outputs_0_aw_valid                ), //o
    .io_outputs_0_aw_ready         (memSub_io_corePorts_0_writeOnly_decoder_io_outputs_0_aw_validPipe_fire), //i
    .io_outputs_0_aw_payload_addr  (io_corePorts_0_writeOnly_decoder_io_outputs_0_aw_payload_addr[31:0]   ), //o
    .io_outputs_0_aw_payload_id    (io_corePorts_0_writeOnly_decoder_io_outputs_0_aw_payload_id[3:0]      ), //o
    .io_outputs_0_aw_payload_len   (io_corePorts_0_writeOnly_decoder_io_outputs_0_aw_payload_len[7:0]     ), //o
    .io_outputs_0_aw_payload_size  (io_corePorts_0_writeOnly_decoder_io_outputs_0_aw_payload_size[2:0]    ), //o
    .io_outputs_0_aw_payload_burst (io_corePorts_0_writeOnly_decoder_io_outputs_0_aw_payload_burst[1:0]   ), //o
    .io_outputs_0_w_valid          (io_corePorts_0_writeOnly_decoder_io_outputs_0_w_valid                 ), //o
    .io_outputs_0_w_ready          (ram_io_axi_arbiter_io_writeInputs_0_w_ready                           ), //i
    .io_outputs_0_w_payload_data   (io_corePorts_0_writeOnly_decoder_io_outputs_0_w_payload_data[31:0]    ), //o
    .io_outputs_0_w_payload_strb   (io_corePorts_0_writeOnly_decoder_io_outputs_0_w_payload_strb[3:0]     ), //o
    .io_outputs_0_w_payload_last   (io_corePorts_0_writeOnly_decoder_io_outputs_0_w_payload_last          ), //o
    .io_outputs_0_b_valid          (ram_io_axi_arbiter_io_writeInputs_0_b_valid                           ), //i
    .io_outputs_0_b_ready          (io_corePorts_0_writeOnly_decoder_io_outputs_0_b_ready                 ), //o
    .io_outputs_0_b_payload_id     (io_corePorts_0_writeOnly_decoder_io_outputs_0_b_payload_id[3:0]       ), //i
    .io_outputs_0_b_payload_resp   (ram_io_axi_arbiter_io_writeInputs_0_b_payload_resp[1:0]               ), //i
    .clk                           (clk                                                                   ), //i
    .reset                         (reset                                                                 )  //i
  );
  Axi4ReadOnlyDecoder io_hostPort_readOnly_decoder (
    .io_input_ar_valid             (io_hostPort_readOnly_ar_valid                                     ), //i
    .io_input_ar_ready             (io_hostPort_readOnly_decoder_io_input_ar_ready                    ), //o
    .io_input_ar_payload_addr      (io_hostPort_readOnly_ar_payload_addr[31:0]                        ), //i
    .io_input_ar_payload_id        (io_hostPort_readOnly_ar_payload_id[3:0]                           ), //i
    .io_input_ar_payload_len       (io_hostPort_readOnly_ar_payload_len[7:0]                          ), //i
    .io_input_ar_payload_size      (io_hostPort_readOnly_ar_payload_size[2:0]                         ), //i
    .io_input_ar_payload_burst     (io_hostPort_readOnly_ar_payload_burst[1:0]                        ), //i
    .io_input_r_valid              (io_hostPort_readOnly_decoder_io_input_r_valid                     ), //o
    .io_input_r_ready              (io_hostPort_readOnly_r_ready                                      ), //i
    .io_input_r_payload_data       (io_hostPort_readOnly_decoder_io_input_r_payload_data[31:0]        ), //o
    .io_input_r_payload_id         (io_hostPort_readOnly_decoder_io_input_r_payload_id[3:0]           ), //o
    .io_input_r_payload_resp       (io_hostPort_readOnly_decoder_io_input_r_payload_resp[1:0]         ), //o
    .io_input_r_payload_last       (io_hostPort_readOnly_decoder_io_input_r_payload_last              ), //o
    .io_outputs_0_ar_valid         (io_hostPort_readOnly_decoder_io_outputs_0_ar_valid                ), //o
    .io_outputs_0_ar_ready         (memSub_io_hostPort_readOnly_decoder_io_outputs_0_ar_validPipe_fire), //i
    .io_outputs_0_ar_payload_addr  (io_hostPort_readOnly_decoder_io_outputs_0_ar_payload_addr[31:0]   ), //o
    .io_outputs_0_ar_payload_id    (io_hostPort_readOnly_decoder_io_outputs_0_ar_payload_id[3:0]      ), //o
    .io_outputs_0_ar_payload_len   (io_hostPort_readOnly_decoder_io_outputs_0_ar_payload_len[7:0]     ), //o
    .io_outputs_0_ar_payload_size  (io_hostPort_readOnly_decoder_io_outputs_0_ar_payload_size[2:0]    ), //o
    .io_outputs_0_ar_payload_burst (io_hostPort_readOnly_decoder_io_outputs_0_ar_payload_burst[1:0]   ), //o
    .io_outputs_0_r_valid          (ram_io_axi_arbiter_io_readInputs_1_r_valid                        ), //i
    .io_outputs_0_r_ready          (io_hostPort_readOnly_decoder_io_outputs_0_r_ready                 ), //o
    .io_outputs_0_r_payload_data   (ram_io_axi_arbiter_io_readInputs_1_r_payload_data[31:0]           ), //i
    .io_outputs_0_r_payload_id     (io_hostPort_readOnly_decoder_io_outputs_0_r_payload_id[3:0]       ), //i
    .io_outputs_0_r_payload_resp   (ram_io_axi_arbiter_io_readInputs_1_r_payload_resp[1:0]            ), //i
    .io_outputs_0_r_payload_last   (ram_io_axi_arbiter_io_readInputs_1_r_payload_last                 ), //i
    .clk                           (clk                                                               ), //i
    .reset                         (reset                                                             )  //i
  );
  Axi4WriteOnlyDecoder io_hostPort_writeOnly_decoder (
    .io_input_aw_valid             (io_hostPort_writeOnly_aw_valid                                     ), //i
    .io_input_aw_ready             (io_hostPort_writeOnly_decoder_io_input_aw_ready                    ), //o
    .io_input_aw_payload_addr      (io_hostPort_writeOnly_aw_payload_addr[31:0]                        ), //i
    .io_input_aw_payload_id        (io_hostPort_writeOnly_aw_payload_id[3:0]                           ), //i
    .io_input_aw_payload_len       (io_hostPort_writeOnly_aw_payload_len[7:0]                          ), //i
    .io_input_aw_payload_size      (io_hostPort_writeOnly_aw_payload_size[2:0]                         ), //i
    .io_input_aw_payload_burst     (io_hostPort_writeOnly_aw_payload_burst[1:0]                        ), //i
    .io_input_w_valid              (io_hostPort_writeOnly_w_valid                                      ), //i
    .io_input_w_ready              (io_hostPort_writeOnly_decoder_io_input_w_ready                     ), //o
    .io_input_w_payload_data       (io_hostPort_writeOnly_w_payload_data[31:0]                         ), //i
    .io_input_w_payload_strb       (io_hostPort_writeOnly_w_payload_strb[3:0]                          ), //i
    .io_input_w_payload_last       (io_hostPort_writeOnly_w_payload_last                               ), //i
    .io_input_b_valid              (io_hostPort_writeOnly_decoder_io_input_b_valid                     ), //o
    .io_input_b_ready              (io_hostPort_writeOnly_b_ready                                      ), //i
    .io_input_b_payload_id         (io_hostPort_writeOnly_decoder_io_input_b_payload_id[3:0]           ), //o
    .io_input_b_payload_resp       (io_hostPort_writeOnly_decoder_io_input_b_payload_resp[1:0]         ), //o
    .io_outputs_0_aw_valid         (io_hostPort_writeOnly_decoder_io_outputs_0_aw_valid                ), //o
    .io_outputs_0_aw_ready         (memSub_io_hostPort_writeOnly_decoder_io_outputs_0_aw_validPipe_fire), //i
    .io_outputs_0_aw_payload_addr  (io_hostPort_writeOnly_decoder_io_outputs_0_aw_payload_addr[31:0]   ), //o
    .io_outputs_0_aw_payload_id    (io_hostPort_writeOnly_decoder_io_outputs_0_aw_payload_id[3:0]      ), //o
    .io_outputs_0_aw_payload_len   (io_hostPort_writeOnly_decoder_io_outputs_0_aw_payload_len[7:0]     ), //o
    .io_outputs_0_aw_payload_size  (io_hostPort_writeOnly_decoder_io_outputs_0_aw_payload_size[2:0]    ), //o
    .io_outputs_0_aw_payload_burst (io_hostPort_writeOnly_decoder_io_outputs_0_aw_payload_burst[1:0]   ), //o
    .io_outputs_0_w_valid          (io_hostPort_writeOnly_decoder_io_outputs_0_w_valid                 ), //o
    .io_outputs_0_w_ready          (ram_io_axi_arbiter_io_writeInputs_1_w_ready                        ), //i
    .io_outputs_0_w_payload_data   (io_hostPort_writeOnly_decoder_io_outputs_0_w_payload_data[31:0]    ), //o
    .io_outputs_0_w_payload_strb   (io_hostPort_writeOnly_decoder_io_outputs_0_w_payload_strb[3:0]     ), //o
    .io_outputs_0_w_payload_last   (io_hostPort_writeOnly_decoder_io_outputs_0_w_payload_last          ), //o
    .io_outputs_0_b_valid          (ram_io_axi_arbiter_io_writeInputs_1_b_valid                        ), //i
    .io_outputs_0_b_ready          (io_hostPort_writeOnly_decoder_io_outputs_0_b_ready                 ), //o
    .io_outputs_0_b_payload_id     (io_hostPort_writeOnly_decoder_io_outputs_0_b_payload_id[3:0]       ), //i
    .io_outputs_0_b_payload_resp   (ram_io_axi_arbiter_io_writeInputs_1_b_payload_resp[1:0]            ), //i
    .clk                           (clk                                                                ), //i
    .reset                         (reset                                                              )  //i
  );
  Axi4SharedArbiter ram_io_axi_arbiter (
    .io_readInputs_0_ar_valid          (memSub_io_corePorts_0_readOnly_decoder_io_outputs_0_ar_validPipe_valid              ), //i
    .io_readInputs_0_ar_ready          (ram_io_axi_arbiter_io_readInputs_0_ar_ready                                         ), //o
    .io_readInputs_0_ar_payload_addr   (ram_io_axi_arbiter_io_readInputs_0_ar_payload_addr[15:0]                            ), //i
    .io_readInputs_0_ar_payload_id     (ram_io_axi_arbiter_io_readInputs_0_ar_payload_id[4:0]                               ), //i
    .io_readInputs_0_ar_payload_len    (memSub_io_corePorts_0_readOnly_decoder_io_outputs_0_ar_validPipe_payload_len[7:0]   ), //i
    .io_readInputs_0_ar_payload_size   (memSub_io_corePorts_0_readOnly_decoder_io_outputs_0_ar_validPipe_payload_size[2:0]  ), //i
    .io_readInputs_0_ar_payload_burst  (memSub_io_corePorts_0_readOnly_decoder_io_outputs_0_ar_validPipe_payload_burst[1:0] ), //i
    .io_readInputs_0_r_valid           (ram_io_axi_arbiter_io_readInputs_0_r_valid                                          ), //o
    .io_readInputs_0_r_ready           (io_corePorts_0_readOnly_decoder_io_outputs_0_r_ready                                ), //i
    .io_readInputs_0_r_payload_data    (ram_io_axi_arbiter_io_readInputs_0_r_payload_data[31:0]                             ), //o
    .io_readInputs_0_r_payload_id      (ram_io_axi_arbiter_io_readInputs_0_r_payload_id[4:0]                                ), //o
    .io_readInputs_0_r_payload_resp    (ram_io_axi_arbiter_io_readInputs_0_r_payload_resp[1:0]                              ), //o
    .io_readInputs_0_r_payload_last    (ram_io_axi_arbiter_io_readInputs_0_r_payload_last                                   ), //o
    .io_readInputs_1_ar_valid          (memSub_io_hostPort_readOnly_decoder_io_outputs_0_ar_validPipe_valid                 ), //i
    .io_readInputs_1_ar_ready          (ram_io_axi_arbiter_io_readInputs_1_ar_ready                                         ), //o
    .io_readInputs_1_ar_payload_addr   (ram_io_axi_arbiter_io_readInputs_1_ar_payload_addr[15:0]                            ), //i
    .io_readInputs_1_ar_payload_id     (ram_io_axi_arbiter_io_readInputs_1_ar_payload_id[4:0]                               ), //i
    .io_readInputs_1_ar_payload_len    (memSub_io_hostPort_readOnly_decoder_io_outputs_0_ar_validPipe_payload_len[7:0]      ), //i
    .io_readInputs_1_ar_payload_size   (memSub_io_hostPort_readOnly_decoder_io_outputs_0_ar_validPipe_payload_size[2:0]     ), //i
    .io_readInputs_1_ar_payload_burst  (memSub_io_hostPort_readOnly_decoder_io_outputs_0_ar_validPipe_payload_burst[1:0]    ), //i
    .io_readInputs_1_r_valid           (ram_io_axi_arbiter_io_readInputs_1_r_valid                                          ), //o
    .io_readInputs_1_r_ready           (io_hostPort_readOnly_decoder_io_outputs_0_r_ready                                   ), //i
    .io_readInputs_1_r_payload_data    (ram_io_axi_arbiter_io_readInputs_1_r_payload_data[31:0]                             ), //o
    .io_readInputs_1_r_payload_id      (ram_io_axi_arbiter_io_readInputs_1_r_payload_id[4:0]                                ), //o
    .io_readInputs_1_r_payload_resp    (ram_io_axi_arbiter_io_readInputs_1_r_payload_resp[1:0]                              ), //o
    .io_readInputs_1_r_payload_last    (ram_io_axi_arbiter_io_readInputs_1_r_payload_last                                   ), //o
    .io_writeInputs_0_aw_valid         (memSub_io_corePorts_0_writeOnly_decoder_io_outputs_0_aw_validPipe_valid             ), //i
    .io_writeInputs_0_aw_ready         (ram_io_axi_arbiter_io_writeInputs_0_aw_ready                                        ), //o
    .io_writeInputs_0_aw_payload_addr  (ram_io_axi_arbiter_io_writeInputs_0_aw_payload_addr[15:0]                           ), //i
    .io_writeInputs_0_aw_payload_id    (ram_io_axi_arbiter_io_writeInputs_0_aw_payload_id[4:0]                              ), //i
    .io_writeInputs_0_aw_payload_len   (memSub_io_corePorts_0_writeOnly_decoder_io_outputs_0_aw_validPipe_payload_len[7:0]  ), //i
    .io_writeInputs_0_aw_payload_size  (memSub_io_corePorts_0_writeOnly_decoder_io_outputs_0_aw_validPipe_payload_size[2:0] ), //i
    .io_writeInputs_0_aw_payload_burst (memSub_io_corePorts_0_writeOnly_decoder_io_outputs_0_aw_validPipe_payload_burst[1:0]), //i
    .io_writeInputs_0_w_valid          (io_corePorts_0_writeOnly_decoder_io_outputs_0_w_valid                               ), //i
    .io_writeInputs_0_w_ready          (ram_io_axi_arbiter_io_writeInputs_0_w_ready                                         ), //o
    .io_writeInputs_0_w_payload_data   (io_corePorts_0_writeOnly_decoder_io_outputs_0_w_payload_data[31:0]                  ), //i
    .io_writeInputs_0_w_payload_strb   (io_corePorts_0_writeOnly_decoder_io_outputs_0_w_payload_strb[3:0]                   ), //i
    .io_writeInputs_0_w_payload_last   (io_corePorts_0_writeOnly_decoder_io_outputs_0_w_payload_last                        ), //i
    .io_writeInputs_0_b_valid          (ram_io_axi_arbiter_io_writeInputs_0_b_valid                                         ), //o
    .io_writeInputs_0_b_ready          (io_corePorts_0_writeOnly_decoder_io_outputs_0_b_ready                               ), //i
    .io_writeInputs_0_b_payload_id     (ram_io_axi_arbiter_io_writeInputs_0_b_payload_id[4:0]                               ), //o
    .io_writeInputs_0_b_payload_resp   (ram_io_axi_arbiter_io_writeInputs_0_b_payload_resp[1:0]                             ), //o
    .io_writeInputs_1_aw_valid         (memSub_io_hostPort_writeOnly_decoder_io_outputs_0_aw_validPipe_valid                ), //i
    .io_writeInputs_1_aw_ready         (ram_io_axi_arbiter_io_writeInputs_1_aw_ready                                        ), //o
    .io_writeInputs_1_aw_payload_addr  (ram_io_axi_arbiter_io_writeInputs_1_aw_payload_addr[15:0]                           ), //i
    .io_writeInputs_1_aw_payload_id    (ram_io_axi_arbiter_io_writeInputs_1_aw_payload_id[4:0]                              ), //i
    .io_writeInputs_1_aw_payload_len   (memSub_io_hostPort_writeOnly_decoder_io_outputs_0_aw_validPipe_payload_len[7:0]     ), //i
    .io_writeInputs_1_aw_payload_size  (memSub_io_hostPort_writeOnly_decoder_io_outputs_0_aw_validPipe_payload_size[2:0]    ), //i
    .io_writeInputs_1_aw_payload_burst (memSub_io_hostPort_writeOnly_decoder_io_outputs_0_aw_validPipe_payload_burst[1:0]   ), //i
    .io_writeInputs_1_w_valid          (io_hostPort_writeOnly_decoder_io_outputs_0_w_valid                                  ), //i
    .io_writeInputs_1_w_ready          (ram_io_axi_arbiter_io_writeInputs_1_w_ready                                         ), //o
    .io_writeInputs_1_w_payload_data   (io_hostPort_writeOnly_decoder_io_outputs_0_w_payload_data[31:0]                     ), //i
    .io_writeInputs_1_w_payload_strb   (io_hostPort_writeOnly_decoder_io_outputs_0_w_payload_strb[3:0]                      ), //i
    .io_writeInputs_1_w_payload_last   (io_hostPort_writeOnly_decoder_io_outputs_0_w_payload_last                           ), //i
    .io_writeInputs_1_b_valid          (ram_io_axi_arbiter_io_writeInputs_1_b_valid                                         ), //o
    .io_writeInputs_1_b_ready          (io_hostPort_writeOnly_decoder_io_outputs_0_b_ready                                  ), //i
    .io_writeInputs_1_b_payload_id     (ram_io_axi_arbiter_io_writeInputs_1_b_payload_id[4:0]                               ), //o
    .io_writeInputs_1_b_payload_resp   (ram_io_axi_arbiter_io_writeInputs_1_b_payload_resp[1:0]                             ), //o
    .io_output_arw_valid               (ram_io_axi_arbiter_io_output_arw_valid                                              ), //o
    .io_output_arw_ready               (ram_io_axi_arw_ready                                                                ), //i
    .io_output_arw_payload_addr        (ram_io_axi_arbiter_io_output_arw_payload_addr[15:0]                                 ), //o
    .io_output_arw_payload_id          (ram_io_axi_arbiter_io_output_arw_payload_id[5:0]                                    ), //o
    .io_output_arw_payload_len         (ram_io_axi_arbiter_io_output_arw_payload_len[7:0]                                   ), //o
    .io_output_arw_payload_size        (ram_io_axi_arbiter_io_output_arw_payload_size[2:0]                                  ), //o
    .io_output_arw_payload_burst       (ram_io_axi_arbiter_io_output_arw_payload_burst[1:0]                                 ), //o
    .io_output_arw_payload_write       (ram_io_axi_arbiter_io_output_arw_payload_write                                      ), //o
    .io_output_w_valid                 (ram_io_axi_arbiter_io_output_w_valid                                                ), //o
    .io_output_w_ready                 (ram_io_axi_w_ready                                                                  ), //i
    .io_output_w_payload_data          (ram_io_axi_arbiter_io_output_w_payload_data[31:0]                                   ), //o
    .io_output_w_payload_strb          (ram_io_axi_arbiter_io_output_w_payload_strb[3:0]                                    ), //o
    .io_output_w_payload_last          (ram_io_axi_arbiter_io_output_w_payload_last                                         ), //o
    .io_output_b_valid                 (ram_io_axi_b_valid                                                                  ), //i
    .io_output_b_ready                 (ram_io_axi_arbiter_io_output_b_ready                                                ), //o
    .io_output_b_payload_id            (ram_io_axi_b_payload_id[5:0]                                                        ), //i
    .io_output_b_payload_resp          (ram_io_axi_b_payload_resp[1:0]                                                      ), //i
    .io_output_r_valid                 (ram_io_axi_r_valid                                                                  ), //i
    .io_output_r_ready                 (ram_io_axi_arbiter_io_output_r_ready                                                ), //o
    .io_output_r_payload_data          (ram_io_axi_r_payload_data[31:0]                                                     ), //i
    .io_output_r_payload_id            (ram_io_axi_r_payload_id[5:0]                                                        ), //i
    .io_output_r_payload_resp          (ram_io_axi_r_payload_resp[1:0]                                                      ), //i
    .io_output_r_payload_last          (ram_io_axi_r_payload_last                                                           ), //i
    .clk                               (clk                                                                                 ), //i
    .reset                             (reset                                                                               )  //i
  );
  assign io_corePorts_0_readOnly_ar_valid = io_corePorts_0_ar_valid;
  assign io_corePorts_0_ar_ready = io_corePorts_0_readOnly_ar_ready;
  assign io_corePorts_0_readOnly_ar_payload_addr = io_corePorts_0_ar_payload_addr;
  assign io_corePorts_0_readOnly_ar_payload_id = io_corePorts_0_ar_payload_id;
  assign io_corePorts_0_readOnly_ar_payload_len = io_corePorts_0_ar_payload_len;
  assign io_corePorts_0_readOnly_ar_payload_size = io_corePorts_0_ar_payload_size;
  assign io_corePorts_0_readOnly_ar_payload_burst = io_corePorts_0_ar_payload_burst;
  assign io_corePorts_0_r_valid = io_corePorts_0_readOnly_r_valid;
  assign io_corePorts_0_readOnly_r_ready = io_corePorts_0_r_ready;
  assign io_corePorts_0_r_payload_data = io_corePorts_0_readOnly_r_payload_data;
  assign io_corePorts_0_r_payload_last = io_corePorts_0_readOnly_r_payload_last;
  assign io_corePorts_0_r_payload_id = io_corePorts_0_readOnly_r_payload_id;
  assign io_corePorts_0_r_payload_resp = io_corePorts_0_readOnly_r_payload_resp;
  assign io_corePorts_0_writeOnly_aw_valid = io_corePorts_0_aw_valid;
  assign io_corePorts_0_aw_ready = io_corePorts_0_writeOnly_aw_ready;
  assign io_corePorts_0_writeOnly_aw_payload_addr = io_corePorts_0_aw_payload_addr;
  assign io_corePorts_0_writeOnly_aw_payload_id = io_corePorts_0_aw_payload_id;
  assign io_corePorts_0_writeOnly_aw_payload_len = io_corePorts_0_aw_payload_len;
  assign io_corePorts_0_writeOnly_aw_payload_size = io_corePorts_0_aw_payload_size;
  assign io_corePorts_0_writeOnly_aw_payload_burst = io_corePorts_0_aw_payload_burst;
  assign io_corePorts_0_writeOnly_w_valid = io_corePorts_0_w_valid;
  assign io_corePorts_0_w_ready = io_corePorts_0_writeOnly_w_ready;
  assign io_corePorts_0_writeOnly_w_payload_data = io_corePorts_0_w_payload_data;
  assign io_corePorts_0_writeOnly_w_payload_strb = io_corePorts_0_w_payload_strb;
  assign io_corePorts_0_writeOnly_w_payload_last = io_corePorts_0_w_payload_last;
  assign io_corePorts_0_b_valid = io_corePorts_0_writeOnly_b_valid;
  assign io_corePorts_0_writeOnly_b_ready = io_corePorts_0_b_ready;
  assign io_corePorts_0_b_payload_id = io_corePorts_0_writeOnly_b_payload_id;
  assign io_corePorts_0_b_payload_resp = io_corePorts_0_writeOnly_b_payload_resp;
  assign io_hostPort_readOnly_ar_valid = io_hostPort_ar_valid;
  assign io_hostPort_ar_ready = io_hostPort_readOnly_ar_ready;
  assign io_hostPort_readOnly_ar_payload_addr = io_hostPort_ar_payload_addr;
  assign io_hostPort_readOnly_ar_payload_id = io_hostPort_ar_payload_id;
  assign io_hostPort_readOnly_ar_payload_len = io_hostPort_ar_payload_len;
  assign io_hostPort_readOnly_ar_payload_size = io_hostPort_ar_payload_size;
  assign io_hostPort_readOnly_ar_payload_burst = io_hostPort_ar_payload_burst;
  assign io_hostPort_r_valid = io_hostPort_readOnly_r_valid;
  assign io_hostPort_readOnly_r_ready = io_hostPort_r_ready;
  assign io_hostPort_r_payload_data = io_hostPort_readOnly_r_payload_data;
  assign io_hostPort_r_payload_last = io_hostPort_readOnly_r_payload_last;
  assign io_hostPort_r_payload_id = io_hostPort_readOnly_r_payload_id;
  assign io_hostPort_r_payload_resp = io_hostPort_readOnly_r_payload_resp;
  assign io_hostPort_writeOnly_aw_valid = io_hostPort_aw_valid;
  assign io_hostPort_aw_ready = io_hostPort_writeOnly_aw_ready;
  assign io_hostPort_writeOnly_aw_payload_addr = io_hostPort_aw_payload_addr;
  assign io_hostPort_writeOnly_aw_payload_id = io_hostPort_aw_payload_id;
  assign io_hostPort_writeOnly_aw_payload_len = io_hostPort_aw_payload_len;
  assign io_hostPort_writeOnly_aw_payload_size = io_hostPort_aw_payload_size;
  assign io_hostPort_writeOnly_aw_payload_burst = io_hostPort_aw_payload_burst;
  assign io_hostPort_writeOnly_w_valid = io_hostPort_w_valid;
  assign io_hostPort_w_ready = io_hostPort_writeOnly_w_ready;
  assign io_hostPort_writeOnly_w_payload_data = io_hostPort_w_payload_data;
  assign io_hostPort_writeOnly_w_payload_strb = io_hostPort_w_payload_strb;
  assign io_hostPort_writeOnly_w_payload_last = io_hostPort_w_payload_last;
  assign io_hostPort_b_valid = io_hostPort_writeOnly_b_valid;
  assign io_hostPort_writeOnly_b_ready = io_hostPort_b_ready;
  assign io_hostPort_b_payload_id = io_hostPort_writeOnly_b_payload_id;
  assign io_hostPort_b_payload_resp = io_hostPort_writeOnly_b_payload_resp;
  assign memSub_io_corePorts_0_readOnly_decoder_io_outputs_0_ar_validPipe_fire = (memSub_io_corePorts_0_readOnly_decoder_io_outputs_0_ar_validPipe_valid && memSub_io_corePorts_0_readOnly_decoder_io_outputs_0_ar_validPipe_ready);
  assign memSub_io_corePorts_0_readOnly_decoder_io_outputs_0_ar_validPipe_valid = memSub_io_corePorts_0_readOnly_decoder_io_outputs_0_ar_rValid;
  assign memSub_io_corePorts_0_readOnly_decoder_io_outputs_0_ar_validPipe_payload_addr = io_corePorts_0_readOnly_decoder_io_outputs_0_ar_payload_addr;
  assign memSub_io_corePorts_0_readOnly_decoder_io_outputs_0_ar_validPipe_payload_id = io_corePorts_0_readOnly_decoder_io_outputs_0_ar_payload_id;
  assign memSub_io_corePorts_0_readOnly_decoder_io_outputs_0_ar_validPipe_payload_len = io_corePorts_0_readOnly_decoder_io_outputs_0_ar_payload_len;
  assign memSub_io_corePorts_0_readOnly_decoder_io_outputs_0_ar_validPipe_payload_size = io_corePorts_0_readOnly_decoder_io_outputs_0_ar_payload_size;
  assign memSub_io_corePorts_0_readOnly_decoder_io_outputs_0_ar_validPipe_payload_burst = io_corePorts_0_readOnly_decoder_io_outputs_0_ar_payload_burst;
  assign memSub_io_corePorts_0_readOnly_decoder_io_outputs_0_ar_validPipe_ready = ram_io_axi_arbiter_io_readInputs_0_ar_ready;
  assign io_corePorts_0_readOnly_decoder_io_outputs_0_r_payload_id = ram_io_axi_arbiter_io_readInputs_0_r_payload_id[3:0];
  assign io_corePorts_0_readOnly_ar_ready = io_corePorts_0_readOnly_decoder_io_input_ar_ready;
  assign io_corePorts_0_readOnly_r_valid = io_corePorts_0_readOnly_decoder_io_input_r_valid;
  assign io_corePorts_0_readOnly_r_payload_data = io_corePorts_0_readOnly_decoder_io_input_r_payload_data;
  assign io_corePorts_0_readOnly_r_payload_last = io_corePorts_0_readOnly_decoder_io_input_r_payload_last;
  assign io_corePorts_0_readOnly_r_payload_id = io_corePorts_0_readOnly_decoder_io_input_r_payload_id;
  assign io_corePorts_0_readOnly_r_payload_resp = io_corePorts_0_readOnly_decoder_io_input_r_payload_resp;
  assign memSub_io_corePorts_0_writeOnly_decoder_io_outputs_0_aw_validPipe_fire = (memSub_io_corePorts_0_writeOnly_decoder_io_outputs_0_aw_validPipe_valid && memSub_io_corePorts_0_writeOnly_decoder_io_outputs_0_aw_validPipe_ready);
  assign memSub_io_corePorts_0_writeOnly_decoder_io_outputs_0_aw_validPipe_valid = memSub_io_corePorts_0_writeOnly_decoder_io_outputs_0_aw_rValid;
  assign memSub_io_corePorts_0_writeOnly_decoder_io_outputs_0_aw_validPipe_payload_addr = io_corePorts_0_writeOnly_decoder_io_outputs_0_aw_payload_addr;
  assign memSub_io_corePorts_0_writeOnly_decoder_io_outputs_0_aw_validPipe_payload_id = io_corePorts_0_writeOnly_decoder_io_outputs_0_aw_payload_id;
  assign memSub_io_corePorts_0_writeOnly_decoder_io_outputs_0_aw_validPipe_payload_len = io_corePorts_0_writeOnly_decoder_io_outputs_0_aw_payload_len;
  assign memSub_io_corePorts_0_writeOnly_decoder_io_outputs_0_aw_validPipe_payload_size = io_corePorts_0_writeOnly_decoder_io_outputs_0_aw_payload_size;
  assign memSub_io_corePorts_0_writeOnly_decoder_io_outputs_0_aw_validPipe_payload_burst = io_corePorts_0_writeOnly_decoder_io_outputs_0_aw_payload_burst;
  assign memSub_io_corePorts_0_writeOnly_decoder_io_outputs_0_aw_validPipe_ready = ram_io_axi_arbiter_io_writeInputs_0_aw_ready;
  assign io_corePorts_0_writeOnly_decoder_io_outputs_0_b_payload_id = ram_io_axi_arbiter_io_writeInputs_0_b_payload_id[3:0];
  assign io_corePorts_0_writeOnly_aw_ready = io_corePorts_0_writeOnly_decoder_io_input_aw_ready;
  assign io_corePorts_0_writeOnly_w_ready = io_corePorts_0_writeOnly_decoder_io_input_w_ready;
  assign io_corePorts_0_writeOnly_b_valid = io_corePorts_0_writeOnly_decoder_io_input_b_valid;
  assign io_corePorts_0_writeOnly_b_payload_id = io_corePorts_0_writeOnly_decoder_io_input_b_payload_id;
  assign io_corePorts_0_writeOnly_b_payload_resp = io_corePorts_0_writeOnly_decoder_io_input_b_payload_resp;
  assign memSub_io_hostPort_readOnly_decoder_io_outputs_0_ar_validPipe_fire = (memSub_io_hostPort_readOnly_decoder_io_outputs_0_ar_validPipe_valid && memSub_io_hostPort_readOnly_decoder_io_outputs_0_ar_validPipe_ready);
  assign memSub_io_hostPort_readOnly_decoder_io_outputs_0_ar_validPipe_valid = memSub_io_hostPort_readOnly_decoder_io_outputs_0_ar_rValid;
  assign memSub_io_hostPort_readOnly_decoder_io_outputs_0_ar_validPipe_payload_addr = io_hostPort_readOnly_decoder_io_outputs_0_ar_payload_addr;
  assign memSub_io_hostPort_readOnly_decoder_io_outputs_0_ar_validPipe_payload_id = io_hostPort_readOnly_decoder_io_outputs_0_ar_payload_id;
  assign memSub_io_hostPort_readOnly_decoder_io_outputs_0_ar_validPipe_payload_len = io_hostPort_readOnly_decoder_io_outputs_0_ar_payload_len;
  assign memSub_io_hostPort_readOnly_decoder_io_outputs_0_ar_validPipe_payload_size = io_hostPort_readOnly_decoder_io_outputs_0_ar_payload_size;
  assign memSub_io_hostPort_readOnly_decoder_io_outputs_0_ar_validPipe_payload_burst = io_hostPort_readOnly_decoder_io_outputs_0_ar_payload_burst;
  assign memSub_io_hostPort_readOnly_decoder_io_outputs_0_ar_validPipe_ready = ram_io_axi_arbiter_io_readInputs_1_ar_ready;
  assign io_hostPort_readOnly_decoder_io_outputs_0_r_payload_id = ram_io_axi_arbiter_io_readInputs_1_r_payload_id[3:0];
  assign io_hostPort_readOnly_ar_ready = io_hostPort_readOnly_decoder_io_input_ar_ready;
  assign io_hostPort_readOnly_r_valid = io_hostPort_readOnly_decoder_io_input_r_valid;
  assign io_hostPort_readOnly_r_payload_data = io_hostPort_readOnly_decoder_io_input_r_payload_data;
  assign io_hostPort_readOnly_r_payload_last = io_hostPort_readOnly_decoder_io_input_r_payload_last;
  assign io_hostPort_readOnly_r_payload_id = io_hostPort_readOnly_decoder_io_input_r_payload_id;
  assign io_hostPort_readOnly_r_payload_resp = io_hostPort_readOnly_decoder_io_input_r_payload_resp;
  assign memSub_io_hostPort_writeOnly_decoder_io_outputs_0_aw_validPipe_fire = (memSub_io_hostPort_writeOnly_decoder_io_outputs_0_aw_validPipe_valid && memSub_io_hostPort_writeOnly_decoder_io_outputs_0_aw_validPipe_ready);
  assign memSub_io_hostPort_writeOnly_decoder_io_outputs_0_aw_validPipe_valid = memSub_io_hostPort_writeOnly_decoder_io_outputs_0_aw_rValid;
  assign memSub_io_hostPort_writeOnly_decoder_io_outputs_0_aw_validPipe_payload_addr = io_hostPort_writeOnly_decoder_io_outputs_0_aw_payload_addr;
  assign memSub_io_hostPort_writeOnly_decoder_io_outputs_0_aw_validPipe_payload_id = io_hostPort_writeOnly_decoder_io_outputs_0_aw_payload_id;
  assign memSub_io_hostPort_writeOnly_decoder_io_outputs_0_aw_validPipe_payload_len = io_hostPort_writeOnly_decoder_io_outputs_0_aw_payload_len;
  assign memSub_io_hostPort_writeOnly_decoder_io_outputs_0_aw_validPipe_payload_size = io_hostPort_writeOnly_decoder_io_outputs_0_aw_payload_size;
  assign memSub_io_hostPort_writeOnly_decoder_io_outputs_0_aw_validPipe_payload_burst = io_hostPort_writeOnly_decoder_io_outputs_0_aw_payload_burst;
  assign memSub_io_hostPort_writeOnly_decoder_io_outputs_0_aw_validPipe_ready = ram_io_axi_arbiter_io_writeInputs_1_aw_ready;
  assign io_hostPort_writeOnly_decoder_io_outputs_0_b_payload_id = ram_io_axi_arbiter_io_writeInputs_1_b_payload_id[3:0];
  assign io_hostPort_writeOnly_aw_ready = io_hostPort_writeOnly_decoder_io_input_aw_ready;
  assign io_hostPort_writeOnly_w_ready = io_hostPort_writeOnly_decoder_io_input_w_ready;
  assign io_hostPort_writeOnly_b_valid = io_hostPort_writeOnly_decoder_io_input_b_valid;
  assign io_hostPort_writeOnly_b_payload_id = io_hostPort_writeOnly_decoder_io_input_b_payload_id;
  assign io_hostPort_writeOnly_b_payload_resp = io_hostPort_writeOnly_decoder_io_input_b_payload_resp;
  assign ram_io_axi_arbiter_io_readInputs_0_ar_payload_addr = memSub_io_corePorts_0_readOnly_decoder_io_outputs_0_ar_validPipe_payload_addr[15:0];
  assign ram_io_axi_arbiter_io_readInputs_0_ar_payload_id = {1'd0, memSub_io_corePorts_0_readOnly_decoder_io_outputs_0_ar_validPipe_payload_id};
  assign ram_io_axi_arbiter_io_readInputs_1_ar_payload_addr = memSub_io_hostPort_readOnly_decoder_io_outputs_0_ar_validPipe_payload_addr[15:0];
  assign ram_io_axi_arbiter_io_readInputs_1_ar_payload_id = {1'd0, memSub_io_hostPort_readOnly_decoder_io_outputs_0_ar_validPipe_payload_id};
  assign ram_io_axi_arbiter_io_writeInputs_0_aw_payload_addr = memSub_io_corePorts_0_writeOnly_decoder_io_outputs_0_aw_validPipe_payload_addr[15:0];
  assign ram_io_axi_arbiter_io_writeInputs_0_aw_payload_id = {1'd0, memSub_io_corePorts_0_writeOnly_decoder_io_outputs_0_aw_validPipe_payload_id};
  assign ram_io_axi_arbiter_io_writeInputs_1_aw_payload_addr = memSub_io_hostPort_writeOnly_decoder_io_outputs_0_aw_validPipe_payload_addr[15:0];
  assign ram_io_axi_arbiter_io_writeInputs_1_aw_payload_id = {1'd0, memSub_io_hostPort_writeOnly_decoder_io_outputs_0_aw_validPipe_payload_id};
  always @(posedge clk) begin
    if(reset) begin
      memSub_io_corePorts_0_readOnly_decoder_io_outputs_0_ar_rValid <= 1'b0;
      memSub_io_corePorts_0_writeOnly_decoder_io_outputs_0_aw_rValid <= 1'b0;
      memSub_io_hostPort_readOnly_decoder_io_outputs_0_ar_rValid <= 1'b0;
      memSub_io_hostPort_writeOnly_decoder_io_outputs_0_aw_rValid <= 1'b0;
    end else begin
      if(io_corePorts_0_readOnly_decoder_io_outputs_0_ar_valid) begin
        memSub_io_corePorts_0_readOnly_decoder_io_outputs_0_ar_rValid <= 1'b1;
      end
      if(memSub_io_corePorts_0_readOnly_decoder_io_outputs_0_ar_validPipe_fire) begin
        memSub_io_corePorts_0_readOnly_decoder_io_outputs_0_ar_rValid <= 1'b0;
      end
      if(io_corePorts_0_writeOnly_decoder_io_outputs_0_aw_valid) begin
        memSub_io_corePorts_0_writeOnly_decoder_io_outputs_0_aw_rValid <= 1'b1;
      end
      if(memSub_io_corePorts_0_writeOnly_decoder_io_outputs_0_aw_validPipe_fire) begin
        memSub_io_corePorts_0_writeOnly_decoder_io_outputs_0_aw_rValid <= 1'b0;
      end
      if(io_hostPort_readOnly_decoder_io_outputs_0_ar_valid) begin
        memSub_io_hostPort_readOnly_decoder_io_outputs_0_ar_rValid <= 1'b1;
      end
      if(memSub_io_hostPort_readOnly_decoder_io_outputs_0_ar_validPipe_fire) begin
        memSub_io_hostPort_readOnly_decoder_io_outputs_0_ar_rValid <= 1'b0;
      end
      if(io_hostPort_writeOnly_decoder_io_outputs_0_aw_valid) begin
        memSub_io_hostPort_writeOnly_decoder_io_outputs_0_aw_rValid <= 1'b1;
      end
      if(memSub_io_hostPort_writeOnly_decoder_io_outputs_0_aw_validPipe_fire) begin
        memSub_io_hostPort_writeOnly_decoder_io_outputs_0_aw_rValid <= 1'b0;
      end
    end
  end


endmodule

module VliwCore (
  input  wire          io_imemWrite_valid,
  input  wire [9:0]    io_imemWrite_payload_addr,
  input  wire [255:0]  io_imemWrite_payload_data,
  output wire          io_dmemAxi_aw_valid,
  input  wire          io_dmemAxi_aw_ready,
  output wire [31:0]   io_dmemAxi_aw_payload_addr,
  output wire [3:0]    io_dmemAxi_aw_payload_id,
  output wire [7:0]    io_dmemAxi_aw_payload_len,
  output wire [2:0]    io_dmemAxi_aw_payload_size,
  output wire [1:0]    io_dmemAxi_aw_payload_burst,
  output wire          io_dmemAxi_w_valid,
  input  wire          io_dmemAxi_w_ready,
  output wire [31:0]   io_dmemAxi_w_payload_data,
  output wire [3:0]    io_dmemAxi_w_payload_strb,
  output wire          io_dmemAxi_w_payload_last,
  input  wire          io_dmemAxi_b_valid,
  output wire          io_dmemAxi_b_ready,
  input  wire [3:0]    io_dmemAxi_b_payload_id,
  input  wire [1:0]    io_dmemAxi_b_payload_resp,
  output wire          io_dmemAxi_ar_valid,
  input  wire          io_dmemAxi_ar_ready,
  output wire [31:0]   io_dmemAxi_ar_payload_addr,
  output wire [3:0]    io_dmemAxi_ar_payload_id,
  output wire [7:0]    io_dmemAxi_ar_payload_len,
  output wire [2:0]    io_dmemAxi_ar_payload_size,
  output wire [1:0]    io_dmemAxi_ar_payload_burst,
  input  wire          io_dmemAxi_r_valid,
  output wire          io_dmemAxi_r_ready,
  input  wire [31:0]   io_dmemAxi_r_payload_data,
  input  wire [3:0]    io_dmemAxi_r_payload_id,
  input  wire [1:0]    io_dmemAxi_r_payload_resp,
  input  wire          io_dmemAxi_r_payload_last,
  input  wire          io_start,
  output wire          io_halted,
  output wire          io_running,
  output wire [9:0]    io_pc,
  output wire          io_wawConflict,
  output wire [31:0]   io_cycleCount,
  input  wire          clk,
  input  wire          reset
);

  wire                fetch_io_stall;
  wire       [10:0]   scratch_io_valuReadAddr_0_0;
  wire       [10:0]   scratch_io_valuReadAddr_0_1;
  wire       [10:0]   scratch_io_valuReadAddr_0_2;
  wire       [10:0]   scratch_io_valuReadAddr_0_3;
  wire       [10:0]   scratch_io_valuReadAddr_0_4;
  wire       [10:0]   scratch_io_valuReadAddr_0_5;
  wire       [10:0]   scratch_io_valuReadAddr_0_6;
  wire       [10:0]   scratch_io_valuReadAddr_0_7;
  wire       [10:0]   scratch_io_valuReadAddr_1_0;
  wire       [10:0]   scratch_io_valuReadAddr_1_1;
  wire       [10:0]   scratch_io_valuReadAddr_1_2;
  wire       [10:0]   scratch_io_valuReadAddr_1_3;
  wire       [10:0]   scratch_io_valuReadAddr_1_4;
  wire       [10:0]   scratch_io_valuReadAddr_1_5;
  wire       [10:0]   scratch_io_valuReadAddr_1_6;
  wire       [10:0]   scratch_io_valuReadAddr_1_7;
  wire       [10:0]   scratch_io_scalarReadAddr_7;
  wire                scratch_io_scalarReadEn_5;
  wire                scratch_io_scalarReadEn_6;
  wire                scratch_io_scalarReadEn_7;
  wire       [255:0]  imem_io_fetchData;
  wire       [9:0]    fetch_io_imemAddr;
  wire       [255:0]  fetch_io_exBundle;
  wire                fetch_io_exValid;
  wire       [9:0]    fetch_io_pc;
  wire                fetch_io_running;
  wire                fetch_io_halted;
  wire                decode_io_aluSlots_0_valid;
  wire       [3:0]    decode_io_aluSlots_0_opcode;
  wire       [10:0]   decode_io_aluSlots_0_dest;
  wire       [10:0]   decode_io_aluSlots_0_src1;
  wire       [10:0]   decode_io_aluSlots_0_src2;
  wire                decode_io_valuSlots_0_valid;
  wire       [3:0]    decode_io_valuSlots_0_opcode;
  wire       [10:0]   decode_io_valuSlots_0_destBase;
  wire       [10:0]   decode_io_valuSlots_0_src1Base;
  wire       [10:0]   decode_io_valuSlots_0_src2Base;
  wire       [10:0]   decode_io_valuSlots_0_src3Base;
  wire                decode_io_loadSlots_0_valid;
  wire       [2:0]    decode_io_loadSlots_0_opcode;
  wire       [10:0]   decode_io_loadSlots_0_dest;
  wire       [10:0]   decode_io_loadSlots_0_addrReg;
  wire       [2:0]    decode_io_loadSlots_0_offset;
  wire       [31:0]   decode_io_loadSlots_0_immediate;
  wire                decode_io_storeSlots_0_valid;
  wire       [1:0]    decode_io_storeSlots_0_opcode;
  wire       [10:0]   decode_io_storeSlots_0_addrReg;
  wire       [10:0]   decode_io_storeSlots_0_srcReg;
  wire                decode_io_flowSlot_valid;
  wire       [3:0]    decode_io_flowSlot_opcode;
  wire       [10:0]   decode_io_flowSlot_dest;
  wire       [10:0]   decode_io_flowSlot_operandA;
  wire       [10:0]   decode_io_flowSlot_operandB;
  wire       [9:0]    decode_io_flowSlot_immediate;
  wire       [31:0]   scratch_io_valuReadData_0_0;
  wire       [31:0]   scratch_io_valuReadData_0_1;
  wire       [31:0]   scratch_io_valuReadData_0_2;
  wire       [31:0]   scratch_io_valuReadData_0_3;
  wire       [31:0]   scratch_io_valuReadData_0_4;
  wire       [31:0]   scratch_io_valuReadData_0_5;
  wire       [31:0]   scratch_io_valuReadData_0_6;
  wire       [31:0]   scratch_io_valuReadData_0_7;
  wire       [31:0]   scratch_io_valuReadData_1_0;
  wire       [31:0]   scratch_io_valuReadData_1_1;
  wire       [31:0]   scratch_io_valuReadData_1_2;
  wire       [31:0]   scratch_io_valuReadData_1_3;
  wire       [31:0]   scratch_io_valuReadData_1_4;
  wire       [31:0]   scratch_io_valuReadData_1_5;
  wire       [31:0]   scratch_io_valuReadData_1_6;
  wire       [31:0]   scratch_io_valuReadData_1_7;
  wire       [31:0]   scratch_io_scalarReadData_0;
  wire       [31:0]   scratch_io_scalarReadData_1;
  wire       [31:0]   scratch_io_scalarReadData_2;
  wire       [31:0]   scratch_io_scalarReadData_3;
  wire       [31:0]   scratch_io_scalarReadData_4;
  wire       [31:0]   scratch_io_scalarReadData_5;
  wire       [31:0]   scratch_io_scalarReadData_6;
  wire       [31:0]   scratch_io_scalarReadData_7;
  wire       [31:0]   scratch_io_scalarReadData_8;
  wire                scratch_io_conflict;
  wire                alu_io_writeReqs_0_valid;
  wire       [10:0]   alu_io_writeReqs_0_payload_addr;
  wire       [31:0]   alu_io_writeReqs_0_payload_data;
  wire                valu_io_writeReqs_0_0_valid;
  wire       [10:0]   valu_io_writeReqs_0_0_payload_addr;
  wire       [31:0]   valu_io_writeReqs_0_0_payload_data;
  wire                valu_io_writeReqs_0_1_valid;
  wire       [10:0]   valu_io_writeReqs_0_1_payload_addr;
  wire       [31:0]   valu_io_writeReqs_0_1_payload_data;
  wire                valu_io_writeReqs_0_2_valid;
  wire       [10:0]   valu_io_writeReqs_0_2_payload_addr;
  wire       [31:0]   valu_io_writeReqs_0_2_payload_data;
  wire                valu_io_writeReqs_0_3_valid;
  wire       [10:0]   valu_io_writeReqs_0_3_payload_addr;
  wire       [31:0]   valu_io_writeReqs_0_3_payload_data;
  wire                valu_io_writeReqs_0_4_valid;
  wire       [10:0]   valu_io_writeReqs_0_4_payload_addr;
  wire       [31:0]   valu_io_writeReqs_0_4_payload_data;
  wire                valu_io_writeReqs_0_5_valid;
  wire       [10:0]   valu_io_writeReqs_0_5_payload_addr;
  wire       [31:0]   valu_io_writeReqs_0_5_payload_data;
  wire                valu_io_writeReqs_0_6_valid;
  wire       [10:0]   valu_io_writeReqs_0_6_payload_addr;
  wire       [31:0]   valu_io_writeReqs_0_6_payload_data;
  wire                valu_io_writeReqs_0_7_valid;
  wire       [10:0]   valu_io_writeReqs_0_7_payload_addr;
  wire       [31:0]   valu_io_writeReqs_0_7_payload_data;
  wire                flow_io_scalarWriteReq_valid;
  wire       [10:0]   flow_io_scalarWriteReq_payload_addr;
  wire       [31:0]   flow_io_scalarWriteReq_payload_data;
  wire                flow_io_vectorWriteReqs_0_valid;
  wire       [10:0]   flow_io_vectorWriteReqs_0_payload_addr;
  wire       [31:0]   flow_io_vectorWriteReqs_0_payload_data;
  wire                flow_io_vectorWriteReqs_1_valid;
  wire       [10:0]   flow_io_vectorWriteReqs_1_payload_addr;
  wire       [31:0]   flow_io_vectorWriteReqs_1_payload_data;
  wire                flow_io_vectorWriteReqs_2_valid;
  wire       [10:0]   flow_io_vectorWriteReqs_2_payload_addr;
  wire       [31:0]   flow_io_vectorWriteReqs_2_payload_data;
  wire                flow_io_vectorWriteReqs_3_valid;
  wire       [10:0]   flow_io_vectorWriteReqs_3_payload_addr;
  wire       [31:0]   flow_io_vectorWriteReqs_3_payload_data;
  wire                flow_io_vectorWriteReqs_4_valid;
  wire       [10:0]   flow_io_vectorWriteReqs_4_payload_addr;
  wire       [31:0]   flow_io_vectorWriteReqs_4_payload_data;
  wire                flow_io_vectorWriteReqs_5_valid;
  wire       [10:0]   flow_io_vectorWriteReqs_5_payload_addr;
  wire       [31:0]   flow_io_vectorWriteReqs_5_payload_data;
  wire                flow_io_vectorWriteReqs_6_valid;
  wire       [10:0]   flow_io_vectorWriteReqs_6_payload_addr;
  wire       [31:0]   flow_io_vectorWriteReqs_6_payload_data;
  wire                flow_io_vectorWriteReqs_7_valid;
  wire       [10:0]   flow_io_vectorWriteReqs_7_payload_addr;
  wire       [31:0]   flow_io_vectorWriteReqs_7_payload_data;
  wire                flow_io_jumpTarget_valid;
  wire       [9:0]    flow_io_jumpTarget_payload;
  wire                flow_io_halt;
  wire                mem_io_axiMaster_ar_valid;
  wire       [31:0]   mem_io_axiMaster_ar_payload_addr;
  wire       [3:0]    mem_io_axiMaster_ar_payload_id;
  wire       [7:0]    mem_io_axiMaster_ar_payload_len;
  wire       [2:0]    mem_io_axiMaster_ar_payload_size;
  wire       [1:0]    mem_io_axiMaster_ar_payload_burst;
  wire                mem_io_axiMaster_aw_valid;
  wire       [31:0]   mem_io_axiMaster_aw_payload_addr;
  wire       [3:0]    mem_io_axiMaster_aw_payload_id;
  wire       [7:0]    mem_io_axiMaster_aw_payload_len;
  wire       [2:0]    mem_io_axiMaster_aw_payload_size;
  wire       [1:0]    mem_io_axiMaster_aw_payload_burst;
  wire                mem_io_axiMaster_w_valid;
  wire       [31:0]   mem_io_axiMaster_w_payload_data;
  wire       [3:0]    mem_io_axiMaster_w_payload_strb;
  wire                mem_io_axiMaster_w_payload_last;
  wire                mem_io_axiMaster_r_ready;
  wire                mem_io_axiMaster_b_ready;
  wire                mem_io_loadWriteReqs_0_valid;
  wire       [10:0]   mem_io_loadWriteReqs_0_payload_addr;
  wire       [31:0]   mem_io_loadWriteReqs_0_payload_data;
  wire                mem_io_constWriteReqs_0_valid;
  wire       [10:0]   mem_io_constWriteReqs_0_payload_addr;
  wire       [31:0]   mem_io_constWriteReqs_0_payload_data;
  wire                mem_io_vloadWriteReqs_0_0_valid;
  wire       [10:0]   mem_io_vloadWriteReqs_0_0_payload_addr;
  wire       [31:0]   mem_io_vloadWriteReqs_0_0_payload_data;
  wire                mem_io_vloadWriteReqs_0_1_valid;
  wire       [10:0]   mem_io_vloadWriteReqs_0_1_payload_addr;
  wire       [31:0]   mem_io_vloadWriteReqs_0_1_payload_data;
  wire                mem_io_vloadWriteReqs_0_2_valid;
  wire       [10:0]   mem_io_vloadWriteReqs_0_2_payload_addr;
  wire       [31:0]   mem_io_vloadWriteReqs_0_2_payload_data;
  wire                mem_io_vloadWriteReqs_0_3_valid;
  wire       [10:0]   mem_io_vloadWriteReqs_0_3_payload_addr;
  wire       [31:0]   mem_io_vloadWriteReqs_0_3_payload_data;
  wire                mem_io_vloadWriteReqs_0_4_valid;
  wire       [10:0]   mem_io_vloadWriteReqs_0_4_payload_addr;
  wire       [31:0]   mem_io_vloadWriteReqs_0_4_payload_data;
  wire                mem_io_vloadWriteReqs_0_5_valid;
  wire       [10:0]   mem_io_vloadWriteReqs_0_5_payload_addr;
  wire       [31:0]   mem_io_vloadWriteReqs_0_5_payload_data;
  wire                mem_io_vloadWriteReqs_0_6_valid;
  wire       [10:0]   mem_io_vloadWriteReqs_0_6_payload_addr;
  wire       [31:0]   mem_io_vloadWriteReqs_0_6_payload_data;
  wire                mem_io_vloadWriteReqs_0_7_valid;
  wire       [10:0]   mem_io_vloadWriteReqs_0_7_payload_addr;
  wire       [31:0]   mem_io_vloadWriteReqs_0_7_payload_data;
  wire                mem_io_stall;
  wire       [10:0]   wb_io_scratchWriteAddr_0;
  wire       [10:0]   wb_io_scratchWriteAddr_1;
  wire       [10:0]   wb_io_scratchWriteAddr_2;
  wire       [10:0]   wb_io_scratchWriteAddr_3;
  wire       [10:0]   wb_io_scratchWriteAddr_4;
  wire       [10:0]   wb_io_scratchWriteAddr_5;
  wire       [10:0]   wb_io_scratchWriteAddr_6;
  wire       [10:0]   wb_io_scratchWriteAddr_7;
  wire       [10:0]   wb_io_scratchWriteAddr_8;
  wire       [10:0]   wb_io_scratchWriteAddr_9;
  wire       [10:0]   wb_io_scratchWriteAddr_10;
  wire       [10:0]   wb_io_scratchWriteAddr_11;
  wire       [10:0]   wb_io_scratchWriteAddr_12;
  wire       [10:0]   wb_io_scratchWriteAddr_13;
  wire       [10:0]   wb_io_scratchWriteAddr_14;
  wire       [10:0]   wb_io_scratchWriteAddr_15;
  wire       [10:0]   wb_io_scratchWriteAddr_16;
  wire       [10:0]   wb_io_scratchWriteAddr_17;
  wire       [10:0]   wb_io_scratchWriteAddr_18;
  wire       [10:0]   wb_io_scratchWriteAddr_19;
  wire       [10:0]   wb_io_scratchWriteAddr_20;
  wire       [10:0]   wb_io_scratchWriteAddr_21;
  wire       [10:0]   wb_io_scratchWriteAddr_22;
  wire       [10:0]   wb_io_scratchWriteAddr_23;
  wire       [10:0]   wb_io_scratchWriteAddr_24;
  wire       [10:0]   wb_io_scratchWriteAddr_25;
  wire       [10:0]   wb_io_scratchWriteAddr_26;
  wire       [10:0]   wb_io_scratchWriteAddr_27;
  wire       [31:0]   wb_io_scratchWriteData_0;
  wire       [31:0]   wb_io_scratchWriteData_1;
  wire       [31:0]   wb_io_scratchWriteData_2;
  wire       [31:0]   wb_io_scratchWriteData_3;
  wire       [31:0]   wb_io_scratchWriteData_4;
  wire       [31:0]   wb_io_scratchWriteData_5;
  wire       [31:0]   wb_io_scratchWriteData_6;
  wire       [31:0]   wb_io_scratchWriteData_7;
  wire       [31:0]   wb_io_scratchWriteData_8;
  wire       [31:0]   wb_io_scratchWriteData_9;
  wire       [31:0]   wb_io_scratchWriteData_10;
  wire       [31:0]   wb_io_scratchWriteData_11;
  wire       [31:0]   wb_io_scratchWriteData_12;
  wire       [31:0]   wb_io_scratchWriteData_13;
  wire       [31:0]   wb_io_scratchWriteData_14;
  wire       [31:0]   wb_io_scratchWriteData_15;
  wire       [31:0]   wb_io_scratchWriteData_16;
  wire       [31:0]   wb_io_scratchWriteData_17;
  wire       [31:0]   wb_io_scratchWriteData_18;
  wire       [31:0]   wb_io_scratchWriteData_19;
  wire       [31:0]   wb_io_scratchWriteData_20;
  wire       [31:0]   wb_io_scratchWriteData_21;
  wire       [31:0]   wb_io_scratchWriteData_22;
  wire       [31:0]   wb_io_scratchWriteData_23;
  wire       [31:0]   wb_io_scratchWriteData_24;
  wire       [31:0]   wb_io_scratchWriteData_25;
  wire       [31:0]   wb_io_scratchWriteData_26;
  wire       [31:0]   wb_io_scratchWriteData_27;
  wire                wb_io_scratchWriteEn_0;
  wire                wb_io_scratchWriteEn_1;
  wire                wb_io_scratchWriteEn_2;
  wire                wb_io_scratchWriteEn_3;
  wire                wb_io_scratchWriteEn_4;
  wire                wb_io_scratchWriteEn_5;
  wire                wb_io_scratchWriteEn_6;
  wire                wb_io_scratchWriteEn_7;
  wire                wb_io_scratchWriteEn_8;
  wire                wb_io_scratchWriteEn_9;
  wire                wb_io_scratchWriteEn_10;
  wire                wb_io_scratchWriteEn_11;
  wire                wb_io_scratchWriteEn_12;
  wire                wb_io_scratchWriteEn_13;
  wire                wb_io_scratchWriteEn_14;
  wire                wb_io_scratchWriteEn_15;
  wire                wb_io_scratchWriteEn_16;
  wire                wb_io_scratchWriteEn_17;
  wire                wb_io_scratchWriteEn_18;
  wire                wb_io_scratchWriteEn_19;
  wire                wb_io_scratchWriteEn_20;
  wire                wb_io_scratchWriteEn_21;
  wire                wb_io_scratchWriteEn_22;
  wire                wb_io_scratchWriteEn_23;
  wire                wb_io_scratchWriteEn_24;
  wire                wb_io_scratchWriteEn_25;
  wire                wb_io_scratchWriteEn_26;
  wire                wb_io_scratchWriteEn_27;
  wire                wb_io_wawConflict;
  reg        [31:0]   cycleCounter;
  reg                 exSlotsReg_valid;
  reg                 exSlotsReg_aluSlots_0_valid;
  reg        [3:0]    exSlotsReg_aluSlots_0_opcode;
  reg        [10:0]   exSlotsReg_aluSlots_0_dest;
  reg        [10:0]   exSlotsReg_aluSlots_0_src1;
  reg        [10:0]   exSlotsReg_aluSlots_0_src2;
  reg                 exSlotsReg_valuSlots_0_valid;
  reg        [3:0]    exSlotsReg_valuSlots_0_opcode;
  reg        [10:0]   exSlotsReg_valuSlots_0_destBase;
  reg        [10:0]   exSlotsReg_valuSlots_0_src1Base;
  reg        [10:0]   exSlotsReg_valuSlots_0_src2Base;
  reg        [10:0]   exSlotsReg_valuSlots_0_src3Base;
  reg                 exSlotsReg_loadSlots_0_valid;
  reg        [2:0]    exSlotsReg_loadSlots_0_opcode;
  reg        [10:0]   exSlotsReg_loadSlots_0_dest;
  reg        [10:0]   exSlotsReg_loadSlots_0_addrReg;
  reg        [2:0]    exSlotsReg_loadSlots_0_offset;
  reg        [31:0]   exSlotsReg_loadSlots_0_immediate;
  reg                 exSlotsReg_storeSlots_0_valid;
  reg        [1:0]    exSlotsReg_storeSlots_0_opcode;
  reg        [10:0]   exSlotsReg_storeSlots_0_addrReg;
  reg        [10:0]   exSlotsReg_storeSlots_0_srcReg;
  reg                 exSlotsReg_flowSlot_valid;
  reg        [3:0]    exSlotsReg_flowSlot_opcode;
  reg        [10:0]   exSlotsReg_flowSlot_dest;
  reg        [10:0]   exSlotsReg_flowSlot_operandA;
  reg        [10:0]   exSlotsReg_flowSlot_operandB;
  reg        [9:0]    exSlotsReg_flowSlot_immediate;
  reg        [9:0]    exSlotsReg_pc;

  InstructionMemory imem (
    .io_fetchAddr          (fetch_io_imemAddr[9:0]          ), //i
    .io_fetchData          (imem_io_fetchData[255:0]        ), //o
    .io_write_valid        (io_imemWrite_valid              ), //i
    .io_write_payload_addr (io_imemWrite_payload_addr[9:0]  ), //i
    .io_write_payload_data (io_imemWrite_payload_data[255:0]), //i
    .clk                   (clk                             ), //i
    .reset                 (reset                           )  //i
  );
  FetchUnit fetch (
    .io_imemAddr     (fetch_io_imemAddr[9:0]         ), //o
    .io_imemData     (imem_io_fetchData[255:0]       ), //i
    .io_exBundle     (fetch_io_exBundle[255:0]       ), //o
    .io_exValid      (fetch_io_exValid               ), //o
    .io_jump_valid   (flow_io_jumpTarget_valid       ), //i
    .io_jump_payload (flow_io_jumpTarget_payload[9:0]), //i
    .io_halt         (flow_io_halt                   ), //i
    .io_start        (io_start                       ), //i
    .io_stall        (fetch_io_stall                 ), //i
    .io_pc           (fetch_io_pc[9:0]               ), //o
    .io_running      (fetch_io_running               ), //o
    .io_halted       (fetch_io_halted                ), //o
    .clk             (clk                            ), //i
    .reset           (reset                          )  //i
  );
  DecodeUnit decode (
    .io_bundle                (fetch_io_exBundle[255:0]             ), //i
    .io_valid                 (fetch_io_exValid                     ), //i
    .io_aluSlots_0_valid      (decode_io_aluSlots_0_valid           ), //o
    .io_aluSlots_0_opcode     (decode_io_aluSlots_0_opcode[3:0]     ), //o
    .io_aluSlots_0_dest       (decode_io_aluSlots_0_dest[10:0]      ), //o
    .io_aluSlots_0_src1       (decode_io_aluSlots_0_src1[10:0]      ), //o
    .io_aluSlots_0_src2       (decode_io_aluSlots_0_src2[10:0]      ), //o
    .io_valuSlots_0_valid     (decode_io_valuSlots_0_valid          ), //o
    .io_valuSlots_0_opcode    (decode_io_valuSlots_0_opcode[3:0]    ), //o
    .io_valuSlots_0_destBase  (decode_io_valuSlots_0_destBase[10:0] ), //o
    .io_valuSlots_0_src1Base  (decode_io_valuSlots_0_src1Base[10:0] ), //o
    .io_valuSlots_0_src2Base  (decode_io_valuSlots_0_src2Base[10:0] ), //o
    .io_valuSlots_0_src3Base  (decode_io_valuSlots_0_src3Base[10:0] ), //o
    .io_loadSlots_0_valid     (decode_io_loadSlots_0_valid          ), //o
    .io_loadSlots_0_opcode    (decode_io_loadSlots_0_opcode[2:0]    ), //o
    .io_loadSlots_0_dest      (decode_io_loadSlots_0_dest[10:0]     ), //o
    .io_loadSlots_0_addrReg   (decode_io_loadSlots_0_addrReg[10:0]  ), //o
    .io_loadSlots_0_offset    (decode_io_loadSlots_0_offset[2:0]    ), //o
    .io_loadSlots_0_immediate (decode_io_loadSlots_0_immediate[31:0]), //o
    .io_storeSlots_0_valid    (decode_io_storeSlots_0_valid         ), //o
    .io_storeSlots_0_opcode   (decode_io_storeSlots_0_opcode[1:0]   ), //o
    .io_storeSlots_0_addrReg  (decode_io_storeSlots_0_addrReg[10:0] ), //o
    .io_storeSlots_0_srcReg   (decode_io_storeSlots_0_srcReg[10:0]  ), //o
    .io_flowSlot_valid        (decode_io_flowSlot_valid             ), //o
    .io_flowSlot_opcode       (decode_io_flowSlot_opcode[3:0]       ), //o
    .io_flowSlot_dest         (decode_io_flowSlot_dest[10:0]        ), //o
    .io_flowSlot_operandA     (decode_io_flowSlot_operandA[10:0]    ), //o
    .io_flowSlot_operandB     (decode_io_flowSlot_operandB[10:0]    ), //o
    .io_flowSlot_immediate    (decode_io_flowSlot_immediate[9:0]    )  //o
  );
  BankedScratchMemory scratch (
    .io_valuReadAddr_0_0 (scratch_io_valuReadAddr_0_0[10:0]   ), //i
    .io_valuReadAddr_0_1 (scratch_io_valuReadAddr_0_1[10:0]   ), //i
    .io_valuReadAddr_0_2 (scratch_io_valuReadAddr_0_2[10:0]   ), //i
    .io_valuReadAddr_0_3 (scratch_io_valuReadAddr_0_3[10:0]   ), //i
    .io_valuReadAddr_0_4 (scratch_io_valuReadAddr_0_4[10:0]   ), //i
    .io_valuReadAddr_0_5 (scratch_io_valuReadAddr_0_5[10:0]   ), //i
    .io_valuReadAddr_0_6 (scratch_io_valuReadAddr_0_6[10:0]   ), //i
    .io_valuReadAddr_0_7 (scratch_io_valuReadAddr_0_7[10:0]   ), //i
    .io_valuReadAddr_1_0 (scratch_io_valuReadAddr_1_0[10:0]   ), //i
    .io_valuReadAddr_1_1 (scratch_io_valuReadAddr_1_1[10:0]   ), //i
    .io_valuReadAddr_1_2 (scratch_io_valuReadAddr_1_2[10:0]   ), //i
    .io_valuReadAddr_1_3 (scratch_io_valuReadAddr_1_3[10:0]   ), //i
    .io_valuReadAddr_1_4 (scratch_io_valuReadAddr_1_4[10:0]   ), //i
    .io_valuReadAddr_1_5 (scratch_io_valuReadAddr_1_5[10:0]   ), //i
    .io_valuReadAddr_1_6 (scratch_io_valuReadAddr_1_6[10:0]   ), //i
    .io_valuReadAddr_1_7 (scratch_io_valuReadAddr_1_7[10:0]   ), //i
    .io_valuReadEn_0_0   (decode_io_valuSlots_0_valid         ), //i
    .io_valuReadEn_0_1   (decode_io_valuSlots_0_valid         ), //i
    .io_valuReadEn_0_2   (decode_io_valuSlots_0_valid         ), //i
    .io_valuReadEn_0_3   (decode_io_valuSlots_0_valid         ), //i
    .io_valuReadEn_0_4   (decode_io_valuSlots_0_valid         ), //i
    .io_valuReadEn_0_5   (decode_io_valuSlots_0_valid         ), //i
    .io_valuReadEn_0_6   (decode_io_valuSlots_0_valid         ), //i
    .io_valuReadEn_0_7   (decode_io_valuSlots_0_valid         ), //i
    .io_valuReadEn_1_0   (decode_io_valuSlots_0_valid         ), //i
    .io_valuReadEn_1_1   (decode_io_valuSlots_0_valid         ), //i
    .io_valuReadEn_1_2   (decode_io_valuSlots_0_valid         ), //i
    .io_valuReadEn_1_3   (decode_io_valuSlots_0_valid         ), //i
    .io_valuReadEn_1_4   (decode_io_valuSlots_0_valid         ), //i
    .io_valuReadEn_1_5   (decode_io_valuSlots_0_valid         ), //i
    .io_valuReadEn_1_6   (decode_io_valuSlots_0_valid         ), //i
    .io_valuReadEn_1_7   (decode_io_valuSlots_0_valid         ), //i
    .io_valuReadData_0_0 (scratch_io_valuReadData_0_0[31:0]   ), //o
    .io_valuReadData_0_1 (scratch_io_valuReadData_0_1[31:0]   ), //o
    .io_valuReadData_0_2 (scratch_io_valuReadData_0_2[31:0]   ), //o
    .io_valuReadData_0_3 (scratch_io_valuReadData_0_3[31:0]   ), //o
    .io_valuReadData_0_4 (scratch_io_valuReadData_0_4[31:0]   ), //o
    .io_valuReadData_0_5 (scratch_io_valuReadData_0_5[31:0]   ), //o
    .io_valuReadData_0_6 (scratch_io_valuReadData_0_6[31:0]   ), //o
    .io_valuReadData_0_7 (scratch_io_valuReadData_0_7[31:0]   ), //o
    .io_valuReadData_1_0 (scratch_io_valuReadData_1_0[31:0]   ), //o
    .io_valuReadData_1_1 (scratch_io_valuReadData_1_1[31:0]   ), //o
    .io_valuReadData_1_2 (scratch_io_valuReadData_1_2[31:0]   ), //o
    .io_valuReadData_1_3 (scratch_io_valuReadData_1_3[31:0]   ), //o
    .io_valuReadData_1_4 (scratch_io_valuReadData_1_4[31:0]   ), //o
    .io_valuReadData_1_5 (scratch_io_valuReadData_1_5[31:0]   ), //o
    .io_valuReadData_1_6 (scratch_io_valuReadData_1_6[31:0]   ), //o
    .io_valuReadData_1_7 (scratch_io_valuReadData_1_7[31:0]   ), //o
    .io_scalarReadAddr_0 (decode_io_aluSlots_0_src1[10:0]     ), //i
    .io_scalarReadAddr_1 (decode_io_aluSlots_0_src2[10:0]     ), //i
    .io_scalarReadAddr_2 (decode_io_loadSlots_0_addrReg[10:0] ), //i
    .io_scalarReadAddr_3 (decode_io_storeSlots_0_addrReg[10:0]), //i
    .io_scalarReadAddr_4 (decode_io_storeSlots_0_srcReg[10:0] ), //i
    .io_scalarReadAddr_5 (decode_io_flowSlot_operandA[10:0]   ), //i
    .io_scalarReadAddr_6 (decode_io_flowSlot_operandB[10:0]   ), //i
    .io_scalarReadAddr_7 (scratch_io_scalarReadAddr_7[10:0]   ), //i
    .io_scalarReadAddr_8 (decode_io_valuSlots_0_src3Base[10:0]), //i
    .io_scalarReadEn_0   (decode_io_aluSlots_0_valid          ), //i
    .io_scalarReadEn_1   (decode_io_aluSlots_0_valid          ), //i
    .io_scalarReadEn_2   (decode_io_loadSlots_0_valid         ), //i
    .io_scalarReadEn_3   (decode_io_storeSlots_0_valid        ), //i
    .io_scalarReadEn_4   (decode_io_storeSlots_0_valid        ), //i
    .io_scalarReadEn_5   (scratch_io_scalarReadEn_5           ), //i
    .io_scalarReadEn_6   (scratch_io_scalarReadEn_6           ), //i
    .io_scalarReadEn_7   (scratch_io_scalarReadEn_7           ), //i
    .io_scalarReadEn_8   (decode_io_valuSlots_0_valid         ), //i
    .io_scalarReadData_0 (scratch_io_scalarReadData_0[31:0]   ), //o
    .io_scalarReadData_1 (scratch_io_scalarReadData_1[31:0]   ), //o
    .io_scalarReadData_2 (scratch_io_scalarReadData_2[31:0]   ), //o
    .io_scalarReadData_3 (scratch_io_scalarReadData_3[31:0]   ), //o
    .io_scalarReadData_4 (scratch_io_scalarReadData_4[31:0]   ), //o
    .io_scalarReadData_5 (scratch_io_scalarReadData_5[31:0]   ), //o
    .io_scalarReadData_6 (scratch_io_scalarReadData_6[31:0]   ), //o
    .io_scalarReadData_7 (scratch_io_scalarReadData_7[31:0]   ), //o
    .io_scalarReadData_8 (scratch_io_scalarReadData_8[31:0]   ), //o
    .io_writeAddr_0      (wb_io_scratchWriteAddr_0[10:0]      ), //i
    .io_writeAddr_1      (wb_io_scratchWriteAddr_1[10:0]      ), //i
    .io_writeAddr_2      (wb_io_scratchWriteAddr_2[10:0]      ), //i
    .io_writeAddr_3      (wb_io_scratchWriteAddr_3[10:0]      ), //i
    .io_writeAddr_4      (wb_io_scratchWriteAddr_4[10:0]      ), //i
    .io_writeAddr_5      (wb_io_scratchWriteAddr_5[10:0]      ), //i
    .io_writeAddr_6      (wb_io_scratchWriteAddr_6[10:0]      ), //i
    .io_writeAddr_7      (wb_io_scratchWriteAddr_7[10:0]      ), //i
    .io_writeAddr_8      (wb_io_scratchWriteAddr_8[10:0]      ), //i
    .io_writeAddr_9      (wb_io_scratchWriteAddr_9[10:0]      ), //i
    .io_writeAddr_10     (wb_io_scratchWriteAddr_10[10:0]     ), //i
    .io_writeAddr_11     (wb_io_scratchWriteAddr_11[10:0]     ), //i
    .io_writeAddr_12     (wb_io_scratchWriteAddr_12[10:0]     ), //i
    .io_writeAddr_13     (wb_io_scratchWriteAddr_13[10:0]     ), //i
    .io_writeAddr_14     (wb_io_scratchWriteAddr_14[10:0]     ), //i
    .io_writeAddr_15     (wb_io_scratchWriteAddr_15[10:0]     ), //i
    .io_writeAddr_16     (wb_io_scratchWriteAddr_16[10:0]     ), //i
    .io_writeAddr_17     (wb_io_scratchWriteAddr_17[10:0]     ), //i
    .io_writeAddr_18     (wb_io_scratchWriteAddr_18[10:0]     ), //i
    .io_writeAddr_19     (wb_io_scratchWriteAddr_19[10:0]     ), //i
    .io_writeAddr_20     (wb_io_scratchWriteAddr_20[10:0]     ), //i
    .io_writeAddr_21     (wb_io_scratchWriteAddr_21[10:0]     ), //i
    .io_writeAddr_22     (wb_io_scratchWriteAddr_22[10:0]     ), //i
    .io_writeAddr_23     (wb_io_scratchWriteAddr_23[10:0]     ), //i
    .io_writeAddr_24     (wb_io_scratchWriteAddr_24[10:0]     ), //i
    .io_writeAddr_25     (wb_io_scratchWriteAddr_25[10:0]     ), //i
    .io_writeAddr_26     (wb_io_scratchWriteAddr_26[10:0]     ), //i
    .io_writeAddr_27     (wb_io_scratchWriteAddr_27[10:0]     ), //i
    .io_writeData_0      (wb_io_scratchWriteData_0[31:0]      ), //i
    .io_writeData_1      (wb_io_scratchWriteData_1[31:0]      ), //i
    .io_writeData_2      (wb_io_scratchWriteData_2[31:0]      ), //i
    .io_writeData_3      (wb_io_scratchWriteData_3[31:0]      ), //i
    .io_writeData_4      (wb_io_scratchWriteData_4[31:0]      ), //i
    .io_writeData_5      (wb_io_scratchWriteData_5[31:0]      ), //i
    .io_writeData_6      (wb_io_scratchWriteData_6[31:0]      ), //i
    .io_writeData_7      (wb_io_scratchWriteData_7[31:0]      ), //i
    .io_writeData_8      (wb_io_scratchWriteData_8[31:0]      ), //i
    .io_writeData_9      (wb_io_scratchWriteData_9[31:0]      ), //i
    .io_writeData_10     (wb_io_scratchWriteData_10[31:0]     ), //i
    .io_writeData_11     (wb_io_scratchWriteData_11[31:0]     ), //i
    .io_writeData_12     (wb_io_scratchWriteData_12[31:0]     ), //i
    .io_writeData_13     (wb_io_scratchWriteData_13[31:0]     ), //i
    .io_writeData_14     (wb_io_scratchWriteData_14[31:0]     ), //i
    .io_writeData_15     (wb_io_scratchWriteData_15[31:0]     ), //i
    .io_writeData_16     (wb_io_scratchWriteData_16[31:0]     ), //i
    .io_writeData_17     (wb_io_scratchWriteData_17[31:0]     ), //i
    .io_writeData_18     (wb_io_scratchWriteData_18[31:0]     ), //i
    .io_writeData_19     (wb_io_scratchWriteData_19[31:0]     ), //i
    .io_writeData_20     (wb_io_scratchWriteData_20[31:0]     ), //i
    .io_writeData_21     (wb_io_scratchWriteData_21[31:0]     ), //i
    .io_writeData_22     (wb_io_scratchWriteData_22[31:0]     ), //i
    .io_writeData_23     (wb_io_scratchWriteData_23[31:0]     ), //i
    .io_writeData_24     (wb_io_scratchWriteData_24[31:0]     ), //i
    .io_writeData_25     (wb_io_scratchWriteData_25[31:0]     ), //i
    .io_writeData_26     (wb_io_scratchWriteData_26[31:0]     ), //i
    .io_writeData_27     (wb_io_scratchWriteData_27[31:0]     ), //i
    .io_writeEn_0        (wb_io_scratchWriteEn_0              ), //i
    .io_writeEn_1        (wb_io_scratchWriteEn_1              ), //i
    .io_writeEn_2        (wb_io_scratchWriteEn_2              ), //i
    .io_writeEn_3        (wb_io_scratchWriteEn_3              ), //i
    .io_writeEn_4        (wb_io_scratchWriteEn_4              ), //i
    .io_writeEn_5        (wb_io_scratchWriteEn_5              ), //i
    .io_writeEn_6        (wb_io_scratchWriteEn_6              ), //i
    .io_writeEn_7        (wb_io_scratchWriteEn_7              ), //i
    .io_writeEn_8        (wb_io_scratchWriteEn_8              ), //i
    .io_writeEn_9        (wb_io_scratchWriteEn_9              ), //i
    .io_writeEn_10       (wb_io_scratchWriteEn_10             ), //i
    .io_writeEn_11       (wb_io_scratchWriteEn_11             ), //i
    .io_writeEn_12       (wb_io_scratchWriteEn_12             ), //i
    .io_writeEn_13       (wb_io_scratchWriteEn_13             ), //i
    .io_writeEn_14       (wb_io_scratchWriteEn_14             ), //i
    .io_writeEn_15       (wb_io_scratchWriteEn_15             ), //i
    .io_writeEn_16       (wb_io_scratchWriteEn_16             ), //i
    .io_writeEn_17       (wb_io_scratchWriteEn_17             ), //i
    .io_writeEn_18       (wb_io_scratchWriteEn_18             ), //i
    .io_writeEn_19       (wb_io_scratchWriteEn_19             ), //i
    .io_writeEn_20       (wb_io_scratchWriteEn_20             ), //i
    .io_writeEn_21       (wb_io_scratchWriteEn_21             ), //i
    .io_writeEn_22       (wb_io_scratchWriteEn_22             ), //i
    .io_writeEn_23       (wb_io_scratchWriteEn_23             ), //i
    .io_writeEn_24       (wb_io_scratchWriteEn_24             ), //i
    .io_writeEn_25       (wb_io_scratchWriteEn_25             ), //i
    .io_writeEn_26       (wb_io_scratchWriteEn_26             ), //i
    .io_writeEn_27       (wb_io_scratchWriteEn_27             ), //i
    .io_conflict         (scratch_io_conflict                 ), //o
    .clk                 (clk                                 ), //i
    .reset               (reset                               )  //i
  );
  AluEngine alu (
    .io_slots_0_valid            (exSlotsReg_aluSlots_0_valid          ), //i
    .io_slots_0_opcode           (exSlotsReg_aluSlots_0_opcode[3:0]    ), //i
    .io_slots_0_dest             (exSlotsReg_aluSlots_0_dest[10:0]     ), //i
    .io_slots_0_src1             (exSlotsReg_aluSlots_0_src1[10:0]     ), //i
    .io_slots_0_src2             (exSlotsReg_aluSlots_0_src2[10:0]     ), //i
    .io_valid                    (exSlotsReg_valid                     ), //i
    .io_operandA_0               (scratch_io_scalarReadData_0[31:0]    ), //i
    .io_operandB_0               (scratch_io_scalarReadData_1[31:0]    ), //i
    .io_writeReqs_0_valid        (alu_io_writeReqs_0_valid             ), //o
    .io_writeReqs_0_payload_addr (alu_io_writeReqs_0_payload_addr[10:0]), //o
    .io_writeReqs_0_payload_data (alu_io_writeReqs_0_payload_data[31:0]), //o
    .clk                         (clk                                  ), //i
    .reset                       (reset                                )  //i
  );
  ValuEngine valu (
    .io_slots_0_valid              (exSlotsReg_valuSlots_0_valid            ), //i
    .io_slots_0_opcode             (exSlotsReg_valuSlots_0_opcode[3:0]      ), //i
    .io_slots_0_destBase           (exSlotsReg_valuSlots_0_destBase[10:0]   ), //i
    .io_slots_0_src1Base           (exSlotsReg_valuSlots_0_src1Base[10:0]   ), //i
    .io_slots_0_src2Base           (exSlotsReg_valuSlots_0_src2Base[10:0]   ), //i
    .io_slots_0_src3Base           (exSlotsReg_valuSlots_0_src3Base[10:0]   ), //i
    .io_valid                      (exSlotsReg_valid                        ), //i
    .io_operandA_0_0               (scratch_io_valuReadData_0_0[31:0]       ), //i
    .io_operandA_0_1               (scratch_io_valuReadData_0_1[31:0]       ), //i
    .io_operandA_0_2               (scratch_io_valuReadData_0_2[31:0]       ), //i
    .io_operandA_0_3               (scratch_io_valuReadData_0_3[31:0]       ), //i
    .io_operandA_0_4               (scratch_io_valuReadData_0_4[31:0]       ), //i
    .io_operandA_0_5               (scratch_io_valuReadData_0_5[31:0]       ), //i
    .io_operandA_0_6               (scratch_io_valuReadData_0_6[31:0]       ), //i
    .io_operandA_0_7               (scratch_io_valuReadData_0_7[31:0]       ), //i
    .io_operandB_0_0               (scratch_io_valuReadData_1_0[31:0]       ), //i
    .io_operandB_0_1               (scratch_io_valuReadData_1_1[31:0]       ), //i
    .io_operandB_0_2               (scratch_io_valuReadData_1_2[31:0]       ), //i
    .io_operandB_0_3               (scratch_io_valuReadData_1_3[31:0]       ), //i
    .io_operandB_0_4               (scratch_io_valuReadData_1_4[31:0]       ), //i
    .io_operandB_0_5               (scratch_io_valuReadData_1_5[31:0]       ), //i
    .io_operandB_0_6               (scratch_io_valuReadData_1_6[31:0]       ), //i
    .io_operandB_0_7               (scratch_io_valuReadData_1_7[31:0]       ), //i
    .io_operandC_0_0               (scratch_io_scalarReadData_8[31:0]       ), //i
    .io_operandC_0_1               (scratch_io_scalarReadData_8[31:0]       ), //i
    .io_operandC_0_2               (scratch_io_scalarReadData_8[31:0]       ), //i
    .io_operandC_0_3               (scratch_io_scalarReadData_8[31:0]       ), //i
    .io_operandC_0_4               (scratch_io_scalarReadData_8[31:0]       ), //i
    .io_operandC_0_5               (scratch_io_scalarReadData_8[31:0]       ), //i
    .io_operandC_0_6               (scratch_io_scalarReadData_8[31:0]       ), //i
    .io_operandC_0_7               (scratch_io_scalarReadData_8[31:0]       ), //i
    .io_writeReqs_0_0_valid        (valu_io_writeReqs_0_0_valid             ), //o
    .io_writeReqs_0_0_payload_addr (valu_io_writeReqs_0_0_payload_addr[10:0]), //o
    .io_writeReqs_0_0_payload_data (valu_io_writeReqs_0_0_payload_data[31:0]), //o
    .io_writeReqs_0_1_valid        (valu_io_writeReqs_0_1_valid             ), //o
    .io_writeReqs_0_1_payload_addr (valu_io_writeReqs_0_1_payload_addr[10:0]), //o
    .io_writeReqs_0_1_payload_data (valu_io_writeReqs_0_1_payload_data[31:0]), //o
    .io_writeReqs_0_2_valid        (valu_io_writeReqs_0_2_valid             ), //o
    .io_writeReqs_0_2_payload_addr (valu_io_writeReqs_0_2_payload_addr[10:0]), //o
    .io_writeReqs_0_2_payload_data (valu_io_writeReqs_0_2_payload_data[31:0]), //o
    .io_writeReqs_0_3_valid        (valu_io_writeReqs_0_3_valid             ), //o
    .io_writeReqs_0_3_payload_addr (valu_io_writeReqs_0_3_payload_addr[10:0]), //o
    .io_writeReqs_0_3_payload_data (valu_io_writeReqs_0_3_payload_data[31:0]), //o
    .io_writeReqs_0_4_valid        (valu_io_writeReqs_0_4_valid             ), //o
    .io_writeReqs_0_4_payload_addr (valu_io_writeReqs_0_4_payload_addr[10:0]), //o
    .io_writeReqs_0_4_payload_data (valu_io_writeReqs_0_4_payload_data[31:0]), //o
    .io_writeReqs_0_5_valid        (valu_io_writeReqs_0_5_valid             ), //o
    .io_writeReqs_0_5_payload_addr (valu_io_writeReqs_0_5_payload_addr[10:0]), //o
    .io_writeReqs_0_5_payload_data (valu_io_writeReqs_0_5_payload_data[31:0]), //o
    .io_writeReqs_0_6_valid        (valu_io_writeReqs_0_6_valid             ), //o
    .io_writeReqs_0_6_payload_addr (valu_io_writeReqs_0_6_payload_addr[10:0]), //o
    .io_writeReqs_0_6_payload_data (valu_io_writeReqs_0_6_payload_data[31:0]), //o
    .io_writeReqs_0_7_valid        (valu_io_writeReqs_0_7_valid             ), //o
    .io_writeReqs_0_7_payload_addr (valu_io_writeReqs_0_7_payload_addr[10:0]), //o
    .io_writeReqs_0_7_payload_data (valu_io_writeReqs_0_7_payload_data[31:0]), //o
    .clk                           (clk                                     ), //i
    .reset                         (reset                                   )  //i
  );
  FlowEngine flow (
    .io_slot_valid                     (exSlotsReg_flowSlot_valid                   ), //i
    .io_slot_opcode                    (exSlotsReg_flowSlot_opcode[3:0]             ), //i
    .io_slot_dest                      (exSlotsReg_flowSlot_dest[10:0]              ), //i
    .io_slot_operandA                  (exSlotsReg_flowSlot_operandA[10:0]          ), //i
    .io_slot_operandB                  (exSlotsReg_flowSlot_operandB[10:0]          ), //i
    .io_slot_immediate                 (exSlotsReg_flowSlot_immediate[9:0]          ), //i
    .io_valid                          (exSlotsReg_valid                            ), //i
    .io_currentPc                      (exSlotsReg_pc[9:0]                          ), //i
    .io_operandCond                    (scratch_io_scalarReadData_5[31:0]           ), //i
    .io_operandA                       (scratch_io_scalarReadData_6[31:0]           ), //i
    .io_operandB                       (scratch_io_scalarReadData_7[31:0]           ), //i
    .io_vCond_0                        (32'h0                                       ), //i
    .io_vCond_1                        (32'h0                                       ), //i
    .io_vCond_2                        (32'h0                                       ), //i
    .io_vCond_3                        (32'h0                                       ), //i
    .io_vCond_4                        (32'h0                                       ), //i
    .io_vCond_5                        (32'h0                                       ), //i
    .io_vCond_6                        (32'h0                                       ), //i
    .io_vCond_7                        (32'h0                                       ), //i
    .io_vSrcA_0                        (32'h0                                       ), //i
    .io_vSrcA_1                        (32'h0                                       ), //i
    .io_vSrcA_2                        (32'h0                                       ), //i
    .io_vSrcA_3                        (32'h0                                       ), //i
    .io_vSrcA_4                        (32'h0                                       ), //i
    .io_vSrcA_5                        (32'h0                                       ), //i
    .io_vSrcA_6                        (32'h0                                       ), //i
    .io_vSrcA_7                        (32'h0                                       ), //i
    .io_vSrcB_0                        (32'h0                                       ), //i
    .io_vSrcB_1                        (32'h0                                       ), //i
    .io_vSrcB_2                        (32'h0                                       ), //i
    .io_vSrcB_3                        (32'h0                                       ), //i
    .io_vSrcB_4                        (32'h0                                       ), //i
    .io_vSrcB_5                        (32'h0                                       ), //i
    .io_vSrcB_6                        (32'h0                                       ), //i
    .io_vSrcB_7                        (32'h0                                       ), //i
    .io_scalarWriteReq_valid           (flow_io_scalarWriteReq_valid                ), //o
    .io_scalarWriteReq_payload_addr    (flow_io_scalarWriteReq_payload_addr[10:0]   ), //o
    .io_scalarWriteReq_payload_data    (flow_io_scalarWriteReq_payload_data[31:0]   ), //o
    .io_vectorWriteReqs_0_valid        (flow_io_vectorWriteReqs_0_valid             ), //o
    .io_vectorWriteReqs_0_payload_addr (flow_io_vectorWriteReqs_0_payload_addr[10:0]), //o
    .io_vectorWriteReqs_0_payload_data (flow_io_vectorWriteReqs_0_payload_data[31:0]), //o
    .io_vectorWriteReqs_1_valid        (flow_io_vectorWriteReqs_1_valid             ), //o
    .io_vectorWriteReqs_1_payload_addr (flow_io_vectorWriteReqs_1_payload_addr[10:0]), //o
    .io_vectorWriteReqs_1_payload_data (flow_io_vectorWriteReqs_1_payload_data[31:0]), //o
    .io_vectorWriteReqs_2_valid        (flow_io_vectorWriteReqs_2_valid             ), //o
    .io_vectorWriteReqs_2_payload_addr (flow_io_vectorWriteReqs_2_payload_addr[10:0]), //o
    .io_vectorWriteReqs_2_payload_data (flow_io_vectorWriteReqs_2_payload_data[31:0]), //o
    .io_vectorWriteReqs_3_valid        (flow_io_vectorWriteReqs_3_valid             ), //o
    .io_vectorWriteReqs_3_payload_addr (flow_io_vectorWriteReqs_3_payload_addr[10:0]), //o
    .io_vectorWriteReqs_3_payload_data (flow_io_vectorWriteReqs_3_payload_data[31:0]), //o
    .io_vectorWriteReqs_4_valid        (flow_io_vectorWriteReqs_4_valid             ), //o
    .io_vectorWriteReqs_4_payload_addr (flow_io_vectorWriteReqs_4_payload_addr[10:0]), //o
    .io_vectorWriteReqs_4_payload_data (flow_io_vectorWriteReqs_4_payload_data[31:0]), //o
    .io_vectorWriteReqs_5_valid        (flow_io_vectorWriteReqs_5_valid             ), //o
    .io_vectorWriteReqs_5_payload_addr (flow_io_vectorWriteReqs_5_payload_addr[10:0]), //o
    .io_vectorWriteReqs_5_payload_data (flow_io_vectorWriteReqs_5_payload_data[31:0]), //o
    .io_vectorWriteReqs_6_valid        (flow_io_vectorWriteReqs_6_valid             ), //o
    .io_vectorWriteReqs_6_payload_addr (flow_io_vectorWriteReqs_6_payload_addr[10:0]), //o
    .io_vectorWriteReqs_6_payload_data (flow_io_vectorWriteReqs_6_payload_data[31:0]), //o
    .io_vectorWriteReqs_7_valid        (flow_io_vectorWriteReqs_7_valid             ), //o
    .io_vectorWriteReqs_7_payload_addr (flow_io_vectorWriteReqs_7_payload_addr[10:0]), //o
    .io_vectorWriteReqs_7_payload_data (flow_io_vectorWriteReqs_7_payload_data[31:0]), //o
    .io_jumpTarget_valid               (flow_io_jumpTarget_valid                    ), //o
    .io_jumpTarget_payload             (flow_io_jumpTarget_payload[9:0]             ), //o
    .io_halt                           (flow_io_halt                                )  //o
  );
  MemoryEngine mem (
    .io_loadSlots_0_valid               (exSlotsReg_loadSlots_0_valid                ), //i
    .io_loadSlots_0_opcode              (exSlotsReg_loadSlots_0_opcode[2:0]          ), //i
    .io_loadSlots_0_dest                (exSlotsReg_loadSlots_0_dest[10:0]           ), //i
    .io_loadSlots_0_addrReg             (exSlotsReg_loadSlots_0_addrReg[10:0]        ), //i
    .io_loadSlots_0_offset              (exSlotsReg_loadSlots_0_offset[2:0]          ), //i
    .io_loadSlots_0_immediate           (exSlotsReg_loadSlots_0_immediate[31:0]      ), //i
    .io_storeSlots_0_valid              (exSlotsReg_storeSlots_0_valid               ), //i
    .io_storeSlots_0_opcode             (exSlotsReg_storeSlots_0_opcode[1:0]         ), //i
    .io_storeSlots_0_addrReg            (exSlotsReg_storeSlots_0_addrReg[10:0]       ), //i
    .io_storeSlots_0_srcReg             (exSlotsReg_storeSlots_0_srcReg[10:0]        ), //i
    .io_valid                           (exSlotsReg_valid                            ), //i
    .io_loadAddrData_0                  (scratch_io_scalarReadData_2[31:0]           ), //i
    .io_storeAddrData_0                 (scratch_io_scalarReadData_3[31:0]           ), //i
    .io_storeSrcData_0                  (scratch_io_scalarReadData_4[31:0]           ), //i
    .io_vstoreSrcData_0_0               (32'h0                                       ), //i
    .io_vstoreSrcData_0_1               (32'h0                                       ), //i
    .io_vstoreSrcData_0_2               (32'h0                                       ), //i
    .io_vstoreSrcData_0_3               (32'h0                                       ), //i
    .io_vstoreSrcData_0_4               (32'h0                                       ), //i
    .io_vstoreSrcData_0_5               (32'h0                                       ), //i
    .io_vstoreSrcData_0_6               (32'h0                                       ), //i
    .io_vstoreSrcData_0_7               (32'h0                                       ), //i
    .io_axiMaster_aw_valid              (mem_io_axiMaster_aw_valid                   ), //o
    .io_axiMaster_aw_ready              (io_dmemAxi_aw_ready                         ), //i
    .io_axiMaster_aw_payload_addr       (mem_io_axiMaster_aw_payload_addr[31:0]      ), //o
    .io_axiMaster_aw_payload_id         (mem_io_axiMaster_aw_payload_id[3:0]         ), //o
    .io_axiMaster_aw_payload_len        (mem_io_axiMaster_aw_payload_len[7:0]        ), //o
    .io_axiMaster_aw_payload_size       (mem_io_axiMaster_aw_payload_size[2:0]       ), //o
    .io_axiMaster_aw_payload_burst      (mem_io_axiMaster_aw_payload_burst[1:0]      ), //o
    .io_axiMaster_w_valid               (mem_io_axiMaster_w_valid                    ), //o
    .io_axiMaster_w_ready               (io_dmemAxi_w_ready                          ), //i
    .io_axiMaster_w_payload_data        (mem_io_axiMaster_w_payload_data[31:0]       ), //o
    .io_axiMaster_w_payload_strb        (mem_io_axiMaster_w_payload_strb[3:0]        ), //o
    .io_axiMaster_w_payload_last        (mem_io_axiMaster_w_payload_last             ), //o
    .io_axiMaster_b_valid               (io_dmemAxi_b_valid                          ), //i
    .io_axiMaster_b_ready               (mem_io_axiMaster_b_ready                    ), //o
    .io_axiMaster_b_payload_id          (io_dmemAxi_b_payload_id[3:0]                ), //i
    .io_axiMaster_b_payload_resp        (io_dmemAxi_b_payload_resp[1:0]              ), //i
    .io_axiMaster_ar_valid              (mem_io_axiMaster_ar_valid                   ), //o
    .io_axiMaster_ar_ready              (io_dmemAxi_ar_ready                         ), //i
    .io_axiMaster_ar_payload_addr       (mem_io_axiMaster_ar_payload_addr[31:0]      ), //o
    .io_axiMaster_ar_payload_id         (mem_io_axiMaster_ar_payload_id[3:0]         ), //o
    .io_axiMaster_ar_payload_len        (mem_io_axiMaster_ar_payload_len[7:0]        ), //o
    .io_axiMaster_ar_payload_size       (mem_io_axiMaster_ar_payload_size[2:0]       ), //o
    .io_axiMaster_ar_payload_burst      (mem_io_axiMaster_ar_payload_burst[1:0]      ), //o
    .io_axiMaster_r_valid               (io_dmemAxi_r_valid                          ), //i
    .io_axiMaster_r_ready               (mem_io_axiMaster_r_ready                    ), //o
    .io_axiMaster_r_payload_data        (io_dmemAxi_r_payload_data[31:0]             ), //i
    .io_axiMaster_r_payload_id          (io_dmemAxi_r_payload_id[3:0]                ), //i
    .io_axiMaster_r_payload_resp        (io_dmemAxi_r_payload_resp[1:0]              ), //i
    .io_axiMaster_r_payload_last        (io_dmemAxi_r_payload_last                   ), //i
    .io_loadWriteReqs_0_valid           (mem_io_loadWriteReqs_0_valid                ), //o
    .io_loadWriteReqs_0_payload_addr    (mem_io_loadWriteReqs_0_payload_addr[10:0]   ), //o
    .io_loadWriteReqs_0_payload_data    (mem_io_loadWriteReqs_0_payload_data[31:0]   ), //o
    .io_constWriteReqs_0_valid          (mem_io_constWriteReqs_0_valid               ), //o
    .io_constWriteReqs_0_payload_addr   (mem_io_constWriteReqs_0_payload_addr[10:0]  ), //o
    .io_constWriteReqs_0_payload_data   (mem_io_constWriteReqs_0_payload_data[31:0]  ), //o
    .io_vloadWriteReqs_0_0_valid        (mem_io_vloadWriteReqs_0_0_valid             ), //o
    .io_vloadWriteReqs_0_0_payload_addr (mem_io_vloadWriteReqs_0_0_payload_addr[10:0]), //o
    .io_vloadWriteReqs_0_0_payload_data (mem_io_vloadWriteReqs_0_0_payload_data[31:0]), //o
    .io_vloadWriteReqs_0_1_valid        (mem_io_vloadWriteReqs_0_1_valid             ), //o
    .io_vloadWriteReqs_0_1_payload_addr (mem_io_vloadWriteReqs_0_1_payload_addr[10:0]), //o
    .io_vloadWriteReqs_0_1_payload_data (mem_io_vloadWriteReqs_0_1_payload_data[31:0]), //o
    .io_vloadWriteReqs_0_2_valid        (mem_io_vloadWriteReqs_0_2_valid             ), //o
    .io_vloadWriteReqs_0_2_payload_addr (mem_io_vloadWriteReqs_0_2_payload_addr[10:0]), //o
    .io_vloadWriteReqs_0_2_payload_data (mem_io_vloadWriteReqs_0_2_payload_data[31:0]), //o
    .io_vloadWriteReqs_0_3_valid        (mem_io_vloadWriteReqs_0_3_valid             ), //o
    .io_vloadWriteReqs_0_3_payload_addr (mem_io_vloadWriteReqs_0_3_payload_addr[10:0]), //o
    .io_vloadWriteReqs_0_3_payload_data (mem_io_vloadWriteReqs_0_3_payload_data[31:0]), //o
    .io_vloadWriteReqs_0_4_valid        (mem_io_vloadWriteReqs_0_4_valid             ), //o
    .io_vloadWriteReqs_0_4_payload_addr (mem_io_vloadWriteReqs_0_4_payload_addr[10:0]), //o
    .io_vloadWriteReqs_0_4_payload_data (mem_io_vloadWriteReqs_0_4_payload_data[31:0]), //o
    .io_vloadWriteReqs_0_5_valid        (mem_io_vloadWriteReqs_0_5_valid             ), //o
    .io_vloadWriteReqs_0_5_payload_addr (mem_io_vloadWriteReqs_0_5_payload_addr[10:0]), //o
    .io_vloadWriteReqs_0_5_payload_data (mem_io_vloadWriteReqs_0_5_payload_data[31:0]), //o
    .io_vloadWriteReqs_0_6_valid        (mem_io_vloadWriteReqs_0_6_valid             ), //o
    .io_vloadWriteReqs_0_6_payload_addr (mem_io_vloadWriteReqs_0_6_payload_addr[10:0]), //o
    .io_vloadWriteReqs_0_6_payload_data (mem_io_vloadWriteReqs_0_6_payload_data[31:0]), //o
    .io_vloadWriteReqs_0_7_valid        (mem_io_vloadWriteReqs_0_7_valid             ), //o
    .io_vloadWriteReqs_0_7_payload_addr (mem_io_vloadWriteReqs_0_7_payload_addr[10:0]), //o
    .io_vloadWriteReqs_0_7_payload_data (mem_io_vloadWriteReqs_0_7_payload_data[31:0]), //o
    .io_stall                           (mem_io_stall                                ), //o
    .clk                                (clk                                         ), //i
    .reset                              (reset                                       )  //i
  );
  WritebackController wb (
    .io_aluWrites_0_valid               (alu_io_writeReqs_0_valid                    ), //i
    .io_aluWrites_0_payload_addr        (alu_io_writeReqs_0_payload_addr[10:0]       ), //i
    .io_aluWrites_0_payload_data        (alu_io_writeReqs_0_payload_data[31:0]       ), //i
    .io_valuWrites_0_valid              (valu_io_writeReqs_0_0_valid                 ), //i
    .io_valuWrites_0_payload_addr       (valu_io_writeReqs_0_0_payload_addr[10:0]    ), //i
    .io_valuWrites_0_payload_data       (valu_io_writeReqs_0_0_payload_data[31:0]    ), //i
    .io_valuWrites_1_valid              (valu_io_writeReqs_0_1_valid                 ), //i
    .io_valuWrites_1_payload_addr       (valu_io_writeReqs_0_1_payload_addr[10:0]    ), //i
    .io_valuWrites_1_payload_data       (valu_io_writeReqs_0_1_payload_data[31:0]    ), //i
    .io_valuWrites_2_valid              (valu_io_writeReqs_0_2_valid                 ), //i
    .io_valuWrites_2_payload_addr       (valu_io_writeReqs_0_2_payload_addr[10:0]    ), //i
    .io_valuWrites_2_payload_data       (valu_io_writeReqs_0_2_payload_data[31:0]    ), //i
    .io_valuWrites_3_valid              (valu_io_writeReqs_0_3_valid                 ), //i
    .io_valuWrites_3_payload_addr       (valu_io_writeReqs_0_3_payload_addr[10:0]    ), //i
    .io_valuWrites_3_payload_data       (valu_io_writeReqs_0_3_payload_data[31:0]    ), //i
    .io_valuWrites_4_valid              (valu_io_writeReqs_0_4_valid                 ), //i
    .io_valuWrites_4_payload_addr       (valu_io_writeReqs_0_4_payload_addr[10:0]    ), //i
    .io_valuWrites_4_payload_data       (valu_io_writeReqs_0_4_payload_data[31:0]    ), //i
    .io_valuWrites_5_valid              (valu_io_writeReqs_0_5_valid                 ), //i
    .io_valuWrites_5_payload_addr       (valu_io_writeReqs_0_5_payload_addr[10:0]    ), //i
    .io_valuWrites_5_payload_data       (valu_io_writeReqs_0_5_payload_data[31:0]    ), //i
    .io_valuWrites_6_valid              (valu_io_writeReqs_0_6_valid                 ), //i
    .io_valuWrites_6_payload_addr       (valu_io_writeReqs_0_6_payload_addr[10:0]    ), //i
    .io_valuWrites_6_payload_data       (valu_io_writeReqs_0_6_payload_data[31:0]    ), //i
    .io_valuWrites_7_valid              (valu_io_writeReqs_0_7_valid                 ), //i
    .io_valuWrites_7_payload_addr       (valu_io_writeReqs_0_7_payload_addr[10:0]    ), //i
    .io_valuWrites_7_payload_data       (valu_io_writeReqs_0_7_payload_data[31:0]    ), //i
    .io_loadWrites_0_valid              (mem_io_loadWriteReqs_0_valid                ), //i
    .io_loadWrites_0_payload_addr       (mem_io_loadWriteReqs_0_payload_addr[10:0]   ), //i
    .io_loadWrites_0_payload_data       (mem_io_loadWriteReqs_0_payload_data[31:0]   ), //i
    .io_constWrites_0_valid             (mem_io_constWriteReqs_0_valid               ), //i
    .io_constWrites_0_payload_addr      (mem_io_constWriteReqs_0_payload_addr[10:0]  ), //i
    .io_constWrites_0_payload_data      (mem_io_constWriteReqs_0_payload_data[31:0]  ), //i
    .io_vloadWrites_0_valid             (mem_io_vloadWriteReqs_0_0_valid             ), //i
    .io_vloadWrites_0_payload_addr      (mem_io_vloadWriteReqs_0_0_payload_addr[10:0]), //i
    .io_vloadWrites_0_payload_data      (mem_io_vloadWriteReqs_0_0_payload_data[31:0]), //i
    .io_vloadWrites_1_valid             (mem_io_vloadWriteReqs_0_1_valid             ), //i
    .io_vloadWrites_1_payload_addr      (mem_io_vloadWriteReqs_0_1_payload_addr[10:0]), //i
    .io_vloadWrites_1_payload_data      (mem_io_vloadWriteReqs_0_1_payload_data[31:0]), //i
    .io_vloadWrites_2_valid             (mem_io_vloadWriteReqs_0_2_valid             ), //i
    .io_vloadWrites_2_payload_addr      (mem_io_vloadWriteReqs_0_2_payload_addr[10:0]), //i
    .io_vloadWrites_2_payload_data      (mem_io_vloadWriteReqs_0_2_payload_data[31:0]), //i
    .io_vloadWrites_3_valid             (mem_io_vloadWriteReqs_0_3_valid             ), //i
    .io_vloadWrites_3_payload_addr      (mem_io_vloadWriteReqs_0_3_payload_addr[10:0]), //i
    .io_vloadWrites_3_payload_data      (mem_io_vloadWriteReqs_0_3_payload_data[31:0]), //i
    .io_vloadWrites_4_valid             (mem_io_vloadWriteReqs_0_4_valid             ), //i
    .io_vloadWrites_4_payload_addr      (mem_io_vloadWriteReqs_0_4_payload_addr[10:0]), //i
    .io_vloadWrites_4_payload_data      (mem_io_vloadWriteReqs_0_4_payload_data[31:0]), //i
    .io_vloadWrites_5_valid             (mem_io_vloadWriteReqs_0_5_valid             ), //i
    .io_vloadWrites_5_payload_addr      (mem_io_vloadWriteReqs_0_5_payload_addr[10:0]), //i
    .io_vloadWrites_5_payload_data      (mem_io_vloadWriteReqs_0_5_payload_data[31:0]), //i
    .io_vloadWrites_6_valid             (mem_io_vloadWriteReqs_0_6_valid             ), //i
    .io_vloadWrites_6_payload_addr      (mem_io_vloadWriteReqs_0_6_payload_addr[10:0]), //i
    .io_vloadWrites_6_payload_data      (mem_io_vloadWriteReqs_0_6_payload_data[31:0]), //i
    .io_vloadWrites_7_valid             (mem_io_vloadWriteReqs_0_7_valid             ), //i
    .io_vloadWrites_7_payload_addr      (mem_io_vloadWriteReqs_0_7_payload_addr[10:0]), //i
    .io_vloadWrites_7_payload_data      (mem_io_vloadWriteReqs_0_7_payload_data[31:0]), //i
    .io_flowScalarWrite_valid           (flow_io_scalarWriteReq_valid                ), //i
    .io_flowScalarWrite_payload_addr    (flow_io_scalarWriteReq_payload_addr[10:0]   ), //i
    .io_flowScalarWrite_payload_data    (flow_io_scalarWriteReq_payload_data[31:0]   ), //i
    .io_flowVectorWrites_0_valid        (flow_io_vectorWriteReqs_0_valid             ), //i
    .io_flowVectorWrites_0_payload_addr (flow_io_vectorWriteReqs_0_payload_addr[10:0]), //i
    .io_flowVectorWrites_0_payload_data (flow_io_vectorWriteReqs_0_payload_data[31:0]), //i
    .io_flowVectorWrites_1_valid        (flow_io_vectorWriteReqs_1_valid             ), //i
    .io_flowVectorWrites_1_payload_addr (flow_io_vectorWriteReqs_1_payload_addr[10:0]), //i
    .io_flowVectorWrites_1_payload_data (flow_io_vectorWriteReqs_1_payload_data[31:0]), //i
    .io_flowVectorWrites_2_valid        (flow_io_vectorWriteReqs_2_valid             ), //i
    .io_flowVectorWrites_2_payload_addr (flow_io_vectorWriteReqs_2_payload_addr[10:0]), //i
    .io_flowVectorWrites_2_payload_data (flow_io_vectorWriteReqs_2_payload_data[31:0]), //i
    .io_flowVectorWrites_3_valid        (flow_io_vectorWriteReqs_3_valid             ), //i
    .io_flowVectorWrites_3_payload_addr (flow_io_vectorWriteReqs_3_payload_addr[10:0]), //i
    .io_flowVectorWrites_3_payload_data (flow_io_vectorWriteReqs_3_payload_data[31:0]), //i
    .io_flowVectorWrites_4_valid        (flow_io_vectorWriteReqs_4_valid             ), //i
    .io_flowVectorWrites_4_payload_addr (flow_io_vectorWriteReqs_4_payload_addr[10:0]), //i
    .io_flowVectorWrites_4_payload_data (flow_io_vectorWriteReqs_4_payload_data[31:0]), //i
    .io_flowVectorWrites_5_valid        (flow_io_vectorWriteReqs_5_valid             ), //i
    .io_flowVectorWrites_5_payload_addr (flow_io_vectorWriteReqs_5_payload_addr[10:0]), //i
    .io_flowVectorWrites_5_payload_data (flow_io_vectorWriteReqs_5_payload_data[31:0]), //i
    .io_flowVectorWrites_6_valid        (flow_io_vectorWriteReqs_6_valid             ), //i
    .io_flowVectorWrites_6_payload_addr (flow_io_vectorWriteReqs_6_payload_addr[10:0]), //i
    .io_flowVectorWrites_6_payload_data (flow_io_vectorWriteReqs_6_payload_data[31:0]), //i
    .io_flowVectorWrites_7_valid        (flow_io_vectorWriteReqs_7_valid             ), //i
    .io_flowVectorWrites_7_payload_addr (flow_io_vectorWriteReqs_7_payload_addr[10:0]), //i
    .io_flowVectorWrites_7_payload_data (flow_io_vectorWriteReqs_7_payload_data[31:0]), //i
    .io_scratchWriteAddr_0              (wb_io_scratchWriteAddr_0[10:0]              ), //o
    .io_scratchWriteAddr_1              (wb_io_scratchWriteAddr_1[10:0]              ), //o
    .io_scratchWriteAddr_2              (wb_io_scratchWriteAddr_2[10:0]              ), //o
    .io_scratchWriteAddr_3              (wb_io_scratchWriteAddr_3[10:0]              ), //o
    .io_scratchWriteAddr_4              (wb_io_scratchWriteAddr_4[10:0]              ), //o
    .io_scratchWriteAddr_5              (wb_io_scratchWriteAddr_5[10:0]              ), //o
    .io_scratchWriteAddr_6              (wb_io_scratchWriteAddr_6[10:0]              ), //o
    .io_scratchWriteAddr_7              (wb_io_scratchWriteAddr_7[10:0]              ), //o
    .io_scratchWriteAddr_8              (wb_io_scratchWriteAddr_8[10:0]              ), //o
    .io_scratchWriteAddr_9              (wb_io_scratchWriteAddr_9[10:0]              ), //o
    .io_scratchWriteAddr_10             (wb_io_scratchWriteAddr_10[10:0]             ), //o
    .io_scratchWriteAddr_11             (wb_io_scratchWriteAddr_11[10:0]             ), //o
    .io_scratchWriteAddr_12             (wb_io_scratchWriteAddr_12[10:0]             ), //o
    .io_scratchWriteAddr_13             (wb_io_scratchWriteAddr_13[10:0]             ), //o
    .io_scratchWriteAddr_14             (wb_io_scratchWriteAddr_14[10:0]             ), //o
    .io_scratchWriteAddr_15             (wb_io_scratchWriteAddr_15[10:0]             ), //o
    .io_scratchWriteAddr_16             (wb_io_scratchWriteAddr_16[10:0]             ), //o
    .io_scratchWriteAddr_17             (wb_io_scratchWriteAddr_17[10:0]             ), //o
    .io_scratchWriteAddr_18             (wb_io_scratchWriteAddr_18[10:0]             ), //o
    .io_scratchWriteAddr_19             (wb_io_scratchWriteAddr_19[10:0]             ), //o
    .io_scratchWriteAddr_20             (wb_io_scratchWriteAddr_20[10:0]             ), //o
    .io_scratchWriteAddr_21             (wb_io_scratchWriteAddr_21[10:0]             ), //o
    .io_scratchWriteAddr_22             (wb_io_scratchWriteAddr_22[10:0]             ), //o
    .io_scratchWriteAddr_23             (wb_io_scratchWriteAddr_23[10:0]             ), //o
    .io_scratchWriteAddr_24             (wb_io_scratchWriteAddr_24[10:0]             ), //o
    .io_scratchWriteAddr_25             (wb_io_scratchWriteAddr_25[10:0]             ), //o
    .io_scratchWriteAddr_26             (wb_io_scratchWriteAddr_26[10:0]             ), //o
    .io_scratchWriteAddr_27             (wb_io_scratchWriteAddr_27[10:0]             ), //o
    .io_scratchWriteData_0              (wb_io_scratchWriteData_0[31:0]              ), //o
    .io_scratchWriteData_1              (wb_io_scratchWriteData_1[31:0]              ), //o
    .io_scratchWriteData_2              (wb_io_scratchWriteData_2[31:0]              ), //o
    .io_scratchWriteData_3              (wb_io_scratchWriteData_3[31:0]              ), //o
    .io_scratchWriteData_4              (wb_io_scratchWriteData_4[31:0]              ), //o
    .io_scratchWriteData_5              (wb_io_scratchWriteData_5[31:0]              ), //o
    .io_scratchWriteData_6              (wb_io_scratchWriteData_6[31:0]              ), //o
    .io_scratchWriteData_7              (wb_io_scratchWriteData_7[31:0]              ), //o
    .io_scratchWriteData_8              (wb_io_scratchWriteData_8[31:0]              ), //o
    .io_scratchWriteData_9              (wb_io_scratchWriteData_9[31:0]              ), //o
    .io_scratchWriteData_10             (wb_io_scratchWriteData_10[31:0]             ), //o
    .io_scratchWriteData_11             (wb_io_scratchWriteData_11[31:0]             ), //o
    .io_scratchWriteData_12             (wb_io_scratchWriteData_12[31:0]             ), //o
    .io_scratchWriteData_13             (wb_io_scratchWriteData_13[31:0]             ), //o
    .io_scratchWriteData_14             (wb_io_scratchWriteData_14[31:0]             ), //o
    .io_scratchWriteData_15             (wb_io_scratchWriteData_15[31:0]             ), //o
    .io_scratchWriteData_16             (wb_io_scratchWriteData_16[31:0]             ), //o
    .io_scratchWriteData_17             (wb_io_scratchWriteData_17[31:0]             ), //o
    .io_scratchWriteData_18             (wb_io_scratchWriteData_18[31:0]             ), //o
    .io_scratchWriteData_19             (wb_io_scratchWriteData_19[31:0]             ), //o
    .io_scratchWriteData_20             (wb_io_scratchWriteData_20[31:0]             ), //o
    .io_scratchWriteData_21             (wb_io_scratchWriteData_21[31:0]             ), //o
    .io_scratchWriteData_22             (wb_io_scratchWriteData_22[31:0]             ), //o
    .io_scratchWriteData_23             (wb_io_scratchWriteData_23[31:0]             ), //o
    .io_scratchWriteData_24             (wb_io_scratchWriteData_24[31:0]             ), //o
    .io_scratchWriteData_25             (wb_io_scratchWriteData_25[31:0]             ), //o
    .io_scratchWriteData_26             (wb_io_scratchWriteData_26[31:0]             ), //o
    .io_scratchWriteData_27             (wb_io_scratchWriteData_27[31:0]             ), //o
    .io_scratchWriteEn_0                (wb_io_scratchWriteEn_0                      ), //o
    .io_scratchWriteEn_1                (wb_io_scratchWriteEn_1                      ), //o
    .io_scratchWriteEn_2                (wb_io_scratchWriteEn_2                      ), //o
    .io_scratchWriteEn_3                (wb_io_scratchWriteEn_3                      ), //o
    .io_scratchWriteEn_4                (wb_io_scratchWriteEn_4                      ), //o
    .io_scratchWriteEn_5                (wb_io_scratchWriteEn_5                      ), //o
    .io_scratchWriteEn_6                (wb_io_scratchWriteEn_6                      ), //o
    .io_scratchWriteEn_7                (wb_io_scratchWriteEn_7                      ), //o
    .io_scratchWriteEn_8                (wb_io_scratchWriteEn_8                      ), //o
    .io_scratchWriteEn_9                (wb_io_scratchWriteEn_9                      ), //o
    .io_scratchWriteEn_10               (wb_io_scratchWriteEn_10                     ), //o
    .io_scratchWriteEn_11               (wb_io_scratchWriteEn_11                     ), //o
    .io_scratchWriteEn_12               (wb_io_scratchWriteEn_12                     ), //o
    .io_scratchWriteEn_13               (wb_io_scratchWriteEn_13                     ), //o
    .io_scratchWriteEn_14               (wb_io_scratchWriteEn_14                     ), //o
    .io_scratchWriteEn_15               (wb_io_scratchWriteEn_15                     ), //o
    .io_scratchWriteEn_16               (wb_io_scratchWriteEn_16                     ), //o
    .io_scratchWriteEn_17               (wb_io_scratchWriteEn_17                     ), //o
    .io_scratchWriteEn_18               (wb_io_scratchWriteEn_18                     ), //o
    .io_scratchWriteEn_19               (wb_io_scratchWriteEn_19                     ), //o
    .io_scratchWriteEn_20               (wb_io_scratchWriteEn_20                     ), //o
    .io_scratchWriteEn_21               (wb_io_scratchWriteEn_21                     ), //o
    .io_scratchWriteEn_22               (wb_io_scratchWriteEn_22                     ), //o
    .io_scratchWriteEn_23               (wb_io_scratchWriteEn_23                     ), //o
    .io_scratchWriteEn_24               (wb_io_scratchWriteEn_24                     ), //o
    .io_scratchWriteEn_25               (wb_io_scratchWriteEn_25                     ), //o
    .io_scratchWriteEn_26               (wb_io_scratchWriteEn_26                     ), //o
    .io_scratchWriteEn_27               (wb_io_scratchWriteEn_27                     ), //o
    .io_wawConflict                     (wb_io_wawConflict                           ), //o
    .clk                                (clk                                         ), //i
    .reset                              (reset                                       )  //i
  );
  assign io_cycleCount = cycleCounter;
  assign scratch_io_scalarReadEn_5 = (decode_io_flowSlot_valid && ((((((decode_io_flowSlot_opcode == 4'b0001) || (decode_io_flowSlot_opcode == 4'b0010)) || (decode_io_flowSlot_opcode == 4'b0011)) || (decode_io_flowSlot_opcode == 4'b0101)) || (decode_io_flowSlot_opcode == 4'b0110)) || (decode_io_flowSlot_opcode == 4'b1000)));
  assign scratch_io_scalarReadEn_6 = (decode_io_flowSlot_valid && ((decode_io_flowSlot_opcode == 4'b0001) || (decode_io_flowSlot_opcode == 4'b0010)));
  assign scratch_io_scalarReadAddr_7 = {1'd0, decode_io_flowSlot_immediate};
  assign scratch_io_scalarReadEn_7 = (decode_io_flowSlot_valid && ((decode_io_flowSlot_opcode == 4'b0001) || (decode_io_flowSlot_opcode == 4'b0010)));
  assign scratch_io_valuReadAddr_0_0 = (decode_io_valuSlots_0_src1Base + 11'h0);
  assign scratch_io_valuReadAddr_0_1 = (decode_io_valuSlots_0_src1Base + 11'h001);
  assign scratch_io_valuReadAddr_0_2 = (decode_io_valuSlots_0_src1Base + 11'h002);
  assign scratch_io_valuReadAddr_0_3 = (decode_io_valuSlots_0_src1Base + 11'h003);
  assign scratch_io_valuReadAddr_0_4 = (decode_io_valuSlots_0_src1Base + 11'h004);
  assign scratch_io_valuReadAddr_0_5 = (decode_io_valuSlots_0_src1Base + 11'h005);
  assign scratch_io_valuReadAddr_0_6 = (decode_io_valuSlots_0_src1Base + 11'h006);
  assign scratch_io_valuReadAddr_0_7 = (decode_io_valuSlots_0_src1Base + 11'h007);
  assign scratch_io_valuReadAddr_1_0 = (decode_io_valuSlots_0_src2Base + 11'h0);
  assign scratch_io_valuReadAddr_1_1 = (decode_io_valuSlots_0_src2Base + 11'h001);
  assign scratch_io_valuReadAddr_1_2 = (decode_io_valuSlots_0_src2Base + 11'h002);
  assign scratch_io_valuReadAddr_1_3 = (decode_io_valuSlots_0_src2Base + 11'h003);
  assign scratch_io_valuReadAddr_1_4 = (decode_io_valuSlots_0_src2Base + 11'h004);
  assign scratch_io_valuReadAddr_1_5 = (decode_io_valuSlots_0_src2Base + 11'h005);
  assign scratch_io_valuReadAddr_1_6 = (decode_io_valuSlots_0_src2Base + 11'h006);
  assign scratch_io_valuReadAddr_1_7 = (decode_io_valuSlots_0_src2Base + 11'h007);
  assign fetch_io_stall = (mem_io_stall || scratch_io_conflict);
  assign io_dmemAxi_aw_valid = mem_io_axiMaster_aw_valid;
  assign io_dmemAxi_aw_payload_addr = mem_io_axiMaster_aw_payload_addr;
  assign io_dmemAxi_aw_payload_id = mem_io_axiMaster_aw_payload_id;
  assign io_dmemAxi_aw_payload_len = mem_io_axiMaster_aw_payload_len;
  assign io_dmemAxi_aw_payload_size = mem_io_axiMaster_aw_payload_size;
  assign io_dmemAxi_aw_payload_burst = mem_io_axiMaster_aw_payload_burst;
  assign io_dmemAxi_w_valid = mem_io_axiMaster_w_valid;
  assign io_dmemAxi_w_payload_data = mem_io_axiMaster_w_payload_data;
  assign io_dmemAxi_w_payload_strb = mem_io_axiMaster_w_payload_strb;
  assign io_dmemAxi_w_payload_last = mem_io_axiMaster_w_payload_last;
  assign io_dmemAxi_b_ready = mem_io_axiMaster_b_ready;
  assign io_dmemAxi_ar_valid = mem_io_axiMaster_ar_valid;
  assign io_dmemAxi_ar_payload_addr = mem_io_axiMaster_ar_payload_addr;
  assign io_dmemAxi_ar_payload_id = mem_io_axiMaster_ar_payload_id;
  assign io_dmemAxi_ar_payload_len = mem_io_axiMaster_ar_payload_len;
  assign io_dmemAxi_ar_payload_size = mem_io_axiMaster_ar_payload_size;
  assign io_dmemAxi_ar_payload_burst = mem_io_axiMaster_ar_payload_burst;
  assign io_dmemAxi_r_ready = mem_io_axiMaster_r_ready;
  assign io_halted = fetch_io_halted;
  assign io_running = fetch_io_running;
  assign io_pc = fetch_io_pc;
  assign io_wawConflict = wb_io_wawConflict;
  always @(posedge clk) begin
    if(reset) begin
      cycleCounter <= 32'h0;
      exSlotsReg_valid <= 1'b0;
      exSlotsReg_pc <= 10'h0;
    end else begin
      if(fetch_io_running) begin
        cycleCounter <= (cycleCounter + 32'h00000001);
      end
      exSlotsReg_valid <= fetch_io_exValid;
      exSlotsReg_pc <= fetch_io_pc;
      if(mem_io_stall) begin
        exSlotsReg_valid <= exSlotsReg_valid;
      end
    end
  end

  always @(posedge clk) begin
    exSlotsReg_aluSlots_0_valid <= decode_io_aluSlots_0_valid;
    exSlotsReg_aluSlots_0_opcode <= decode_io_aluSlots_0_opcode;
    exSlotsReg_aluSlots_0_dest <= decode_io_aluSlots_0_dest;
    exSlotsReg_aluSlots_0_src1 <= decode_io_aluSlots_0_src1;
    exSlotsReg_aluSlots_0_src2 <= decode_io_aluSlots_0_src2;
    exSlotsReg_valuSlots_0_valid <= decode_io_valuSlots_0_valid;
    exSlotsReg_valuSlots_0_opcode <= decode_io_valuSlots_0_opcode;
    exSlotsReg_valuSlots_0_destBase <= decode_io_valuSlots_0_destBase;
    exSlotsReg_valuSlots_0_src1Base <= decode_io_valuSlots_0_src1Base;
    exSlotsReg_valuSlots_0_src2Base <= decode_io_valuSlots_0_src2Base;
    exSlotsReg_valuSlots_0_src3Base <= decode_io_valuSlots_0_src3Base;
    exSlotsReg_loadSlots_0_valid <= decode_io_loadSlots_0_valid;
    exSlotsReg_loadSlots_0_opcode <= decode_io_loadSlots_0_opcode;
    exSlotsReg_loadSlots_0_dest <= decode_io_loadSlots_0_dest;
    exSlotsReg_loadSlots_0_addrReg <= decode_io_loadSlots_0_addrReg;
    exSlotsReg_loadSlots_0_offset <= decode_io_loadSlots_0_offset;
    exSlotsReg_loadSlots_0_immediate <= decode_io_loadSlots_0_immediate;
    exSlotsReg_storeSlots_0_valid <= decode_io_storeSlots_0_valid;
    exSlotsReg_storeSlots_0_opcode <= decode_io_storeSlots_0_opcode;
    exSlotsReg_storeSlots_0_addrReg <= decode_io_storeSlots_0_addrReg;
    exSlotsReg_storeSlots_0_srcReg <= decode_io_storeSlots_0_srcReg;
    exSlotsReg_flowSlot_valid <= decode_io_flowSlot_valid;
    exSlotsReg_flowSlot_opcode <= decode_io_flowSlot_opcode;
    exSlotsReg_flowSlot_dest <= decode_io_flowSlot_dest;
    exSlotsReg_flowSlot_operandA <= decode_io_flowSlot_operandA;
    exSlotsReg_flowSlot_operandB <= decode_io_flowSlot_operandB;
    exSlotsReg_flowSlot_immediate <= decode_io_flowSlot_immediate;
  end


endmodule

module Axi4SharedArbiter (
  input  wire          io_readInputs_0_ar_valid,
  output wire          io_readInputs_0_ar_ready,
  input  wire [15:0]   io_readInputs_0_ar_payload_addr,
  input  wire [4:0]    io_readInputs_0_ar_payload_id,
  input  wire [7:0]    io_readInputs_0_ar_payload_len,
  input  wire [2:0]    io_readInputs_0_ar_payload_size,
  input  wire [1:0]    io_readInputs_0_ar_payload_burst,
  output wire          io_readInputs_0_r_valid,
  input  wire          io_readInputs_0_r_ready,
  output wire [31:0]   io_readInputs_0_r_payload_data,
  output wire [4:0]    io_readInputs_0_r_payload_id,
  output wire [1:0]    io_readInputs_0_r_payload_resp,
  output wire          io_readInputs_0_r_payload_last,
  input  wire          io_readInputs_1_ar_valid,
  output wire          io_readInputs_1_ar_ready,
  input  wire [15:0]   io_readInputs_1_ar_payload_addr,
  input  wire [4:0]    io_readInputs_1_ar_payload_id,
  input  wire [7:0]    io_readInputs_1_ar_payload_len,
  input  wire [2:0]    io_readInputs_1_ar_payload_size,
  input  wire [1:0]    io_readInputs_1_ar_payload_burst,
  output wire          io_readInputs_1_r_valid,
  input  wire          io_readInputs_1_r_ready,
  output wire [31:0]   io_readInputs_1_r_payload_data,
  output wire [4:0]    io_readInputs_1_r_payload_id,
  output wire [1:0]    io_readInputs_1_r_payload_resp,
  output wire          io_readInputs_1_r_payload_last,
  input  wire          io_writeInputs_0_aw_valid,
  output wire          io_writeInputs_0_aw_ready,
  input  wire [15:0]   io_writeInputs_0_aw_payload_addr,
  input  wire [4:0]    io_writeInputs_0_aw_payload_id,
  input  wire [7:0]    io_writeInputs_0_aw_payload_len,
  input  wire [2:0]    io_writeInputs_0_aw_payload_size,
  input  wire [1:0]    io_writeInputs_0_aw_payload_burst,
  input  wire          io_writeInputs_0_w_valid,
  output wire          io_writeInputs_0_w_ready,
  input  wire [31:0]   io_writeInputs_0_w_payload_data,
  input  wire [3:0]    io_writeInputs_0_w_payload_strb,
  input  wire          io_writeInputs_0_w_payload_last,
  output wire          io_writeInputs_0_b_valid,
  input  wire          io_writeInputs_0_b_ready,
  output wire [4:0]    io_writeInputs_0_b_payload_id,
  output wire [1:0]    io_writeInputs_0_b_payload_resp,
  input  wire          io_writeInputs_1_aw_valid,
  output wire          io_writeInputs_1_aw_ready,
  input  wire [15:0]   io_writeInputs_1_aw_payload_addr,
  input  wire [4:0]    io_writeInputs_1_aw_payload_id,
  input  wire [7:0]    io_writeInputs_1_aw_payload_len,
  input  wire [2:0]    io_writeInputs_1_aw_payload_size,
  input  wire [1:0]    io_writeInputs_1_aw_payload_burst,
  input  wire          io_writeInputs_1_w_valid,
  output wire          io_writeInputs_1_w_ready,
  input  wire [31:0]   io_writeInputs_1_w_payload_data,
  input  wire [3:0]    io_writeInputs_1_w_payload_strb,
  input  wire          io_writeInputs_1_w_payload_last,
  output wire          io_writeInputs_1_b_valid,
  input  wire          io_writeInputs_1_b_ready,
  output wire [4:0]    io_writeInputs_1_b_payload_id,
  output wire [1:0]    io_writeInputs_1_b_payload_resp,
  output wire          io_output_arw_valid,
  input  wire          io_output_arw_ready,
  output wire [15:0]   io_output_arw_payload_addr,
  output wire [5:0]    io_output_arw_payload_id,
  output wire [7:0]    io_output_arw_payload_len,
  output wire [2:0]    io_output_arw_payload_size,
  output wire [1:0]    io_output_arw_payload_burst,
  output wire          io_output_arw_payload_write,
  output wire          io_output_w_valid,
  input  wire          io_output_w_ready,
  output wire [31:0]   io_output_w_payload_data,
  output wire [3:0]    io_output_w_payload_strb,
  output wire          io_output_w_payload_last,
  input  wire          io_output_b_valid,
  output wire          io_output_b_ready,
  input  wire [5:0]    io_output_b_payload_id,
  input  wire [1:0]    io_output_b_payload_resp,
  input  wire          io_output_r_valid,
  output wire          io_output_r_ready,
  input  wire [31:0]   io_output_r_payload_data,
  input  wire [5:0]    io_output_r_payload_id,
  input  wire [1:0]    io_output_r_payload_resp,
  input  wire          io_output_r_payload_last,
  input  wire          clk,
  input  wire          reset
);

  reg                 cmdArbiter_io_output_ready;
  wire                cmdRouteFork_thrown_translated_fifo_io_pop_ready;
  wire                cmdArbiter_io_inputs_0_ready;
  wire                cmdArbiter_io_inputs_1_ready;
  wire                cmdArbiter_io_inputs_2_ready;
  wire                cmdArbiter_io_inputs_3_ready;
  wire                cmdArbiter_io_output_valid;
  wire       [15:0]   cmdArbiter_io_output_payload_addr;
  wire       [4:0]    cmdArbiter_io_output_payload_id;
  wire       [7:0]    cmdArbiter_io_output_payload_len;
  wire       [2:0]    cmdArbiter_io_output_payload_size;
  wire       [1:0]    cmdArbiter_io_output_payload_burst;
  wire                cmdArbiter_io_output_payload_write;
  wire       [1:0]    cmdArbiter_io_chosen;
  wire       [3:0]    cmdArbiter_io_chosenOH;
  wire                cmdRouteFork_thrown_translated_fifo_io_push_ready;
  wire                cmdRouteFork_thrown_translated_fifo_io_pop_valid;
  wire       [0:0]    cmdRouteFork_thrown_translated_fifo_io_pop_payload;
  wire       [2:0]    cmdRouteFork_thrown_translated_fifo_io_occupancy;
  wire       [2:0]    cmdRouteFork_thrown_translated_fifo_io_availability;
  wire       [1:0]    _zz__zz_io_output_arw_payload_id;
  wire       [1:0]    _zz__zz_io_output_arw_payload_id_1;
  wire       [1:0]    _zz__zz_cmdRouteFork_thrown_translated_payload;
  reg                 _zz_writeLogic_routeDataInput_valid;
  reg                 _zz_writeLogic_routeDataInput_ready;
  reg        [31:0]   _zz_writeLogic_routeDataInput_payload_data;
  reg        [3:0]    _zz_writeLogic_routeDataInput_payload_strb;
  reg                 _zz_writeLogic_routeDataInput_payload_last;
  reg                 _zz_io_output_b_ready;
  reg                 _zz_io_output_r_ready;
  wire                inputsCmd_0_valid;
  wire                inputsCmd_0_ready;
  wire       [15:0]   inputsCmd_0_payload_addr;
  wire       [4:0]    inputsCmd_0_payload_id;
  wire       [7:0]    inputsCmd_0_payload_len;
  wire       [2:0]    inputsCmd_0_payload_size;
  wire       [1:0]    inputsCmd_0_payload_burst;
  wire                inputsCmd_0_payload_write;
  wire                inputsCmd_1_valid;
  wire                inputsCmd_1_ready;
  wire       [15:0]   inputsCmd_1_payload_addr;
  wire       [4:0]    inputsCmd_1_payload_id;
  wire       [7:0]    inputsCmd_1_payload_len;
  wire       [2:0]    inputsCmd_1_payload_size;
  wire       [1:0]    inputsCmd_1_payload_burst;
  wire                inputsCmd_1_payload_write;
  wire                inputsCmd_2_valid;
  wire                inputsCmd_2_ready;
  wire       [15:0]   inputsCmd_2_payload_addr;
  wire       [4:0]    inputsCmd_2_payload_id;
  wire       [7:0]    inputsCmd_2_payload_len;
  wire       [2:0]    inputsCmd_2_payload_size;
  wire       [1:0]    inputsCmd_2_payload_burst;
  wire                inputsCmd_2_payload_write;
  wire                inputsCmd_3_valid;
  wire                inputsCmd_3_ready;
  wire       [15:0]   inputsCmd_3_payload_addr;
  wire       [4:0]    inputsCmd_3_payload_id;
  wire       [7:0]    inputsCmd_3_payload_len;
  wire       [2:0]    inputsCmd_3_payload_size;
  wire       [1:0]    inputsCmd_3_payload_burst;
  wire                inputsCmd_3_payload_write;
  wire                cmdOutputFork_valid;
  wire                cmdOutputFork_ready;
  wire       [15:0]   cmdOutputFork_payload_addr;
  wire       [4:0]    cmdOutputFork_payload_id;
  wire       [7:0]    cmdOutputFork_payload_len;
  wire       [2:0]    cmdOutputFork_payload_size;
  wire       [1:0]    cmdOutputFork_payload_burst;
  wire                cmdOutputFork_payload_write;
  wire                cmdRouteFork_valid;
  reg                 cmdRouteFork_ready;
  wire       [15:0]   cmdRouteFork_payload_addr;
  wire       [4:0]    cmdRouteFork_payload_id;
  wire       [7:0]    cmdRouteFork_payload_len;
  wire       [2:0]    cmdRouteFork_payload_size;
  wire       [1:0]    cmdRouteFork_payload_burst;
  wire                cmdRouteFork_payload_write;
  reg                 ram_io_axi_arbiter_cmdArbiter_io_output_fork2_logic_linkEnable_0;
  reg                 ram_io_axi_arbiter_cmdArbiter_io_output_fork2_logic_linkEnable_1;
  wire                when_Stream_l1063;
  wire                when_Stream_l1063_1;
  wire                cmdOutputFork_fire;
  wire                cmdRouteFork_fire;
  wire                _zz_io_output_arw_payload_id;
  wire                _zz_io_output_arw_payload_id_1;
  wire                when_Stream_l445;
  reg                 cmdRouteFork_thrown_valid;
  wire                cmdRouteFork_thrown_ready;
  wire       [15:0]   cmdRouteFork_thrown_payload_addr;
  wire       [4:0]    cmdRouteFork_thrown_payload_id;
  wire       [7:0]    cmdRouteFork_thrown_payload_len;
  wire       [2:0]    cmdRouteFork_thrown_payload_size;
  wire       [1:0]    cmdRouteFork_thrown_payload_burst;
  wire                cmdRouteFork_thrown_payload_write;
  wire                _zz_cmdRouteFork_thrown_translated_payload;
  wire                cmdRouteFork_thrown_translated_valid;
  wire                cmdRouteFork_thrown_translated_ready;
  wire       [0:0]    cmdRouteFork_thrown_translated_payload;
  wire                writeLogic_routeDataInput_valid;
  wire                writeLogic_routeDataInput_ready;
  wire       [31:0]   writeLogic_routeDataInput_payload_data;
  wire       [3:0]    writeLogic_routeDataInput_payload_strb;
  wire                writeLogic_routeDataInput_payload_last;
  wire                io_output_w_fire;
  wire       [0:0]    writeLogic_writeRspIndex;
  wire                writeLogic_writeRspSels_0;
  wire                writeLogic_writeRspSels_1;
  wire       [0:0]    readRspIndex;
  wire                readRspSels_0;
  wire                readRspSels_1;

  assign _zz__zz_io_output_arw_payload_id = cmdArbiter_io_chosenOH[3 : 2];
  assign _zz__zz_io_output_arw_payload_id_1 = cmdArbiter_io_chosenOH[1 : 0];
  assign _zz__zz_cmdRouteFork_thrown_translated_payload = cmdArbiter_io_chosenOH[3 : 2];
  StreamArbiter cmdArbiter (
    .io_inputs_0_valid         (inputsCmd_0_valid                      ), //i
    .io_inputs_0_ready         (cmdArbiter_io_inputs_0_ready           ), //o
    .io_inputs_0_payload_addr  (inputsCmd_0_payload_addr[15:0]         ), //i
    .io_inputs_0_payload_id    (inputsCmd_0_payload_id[4:0]            ), //i
    .io_inputs_0_payload_len   (inputsCmd_0_payload_len[7:0]           ), //i
    .io_inputs_0_payload_size  (inputsCmd_0_payload_size[2:0]          ), //i
    .io_inputs_0_payload_burst (inputsCmd_0_payload_burst[1:0]         ), //i
    .io_inputs_0_payload_write (inputsCmd_0_payload_write              ), //i
    .io_inputs_1_valid         (inputsCmd_1_valid                      ), //i
    .io_inputs_1_ready         (cmdArbiter_io_inputs_1_ready           ), //o
    .io_inputs_1_payload_addr  (inputsCmd_1_payload_addr[15:0]         ), //i
    .io_inputs_1_payload_id    (inputsCmd_1_payload_id[4:0]            ), //i
    .io_inputs_1_payload_len   (inputsCmd_1_payload_len[7:0]           ), //i
    .io_inputs_1_payload_size  (inputsCmd_1_payload_size[2:0]          ), //i
    .io_inputs_1_payload_burst (inputsCmd_1_payload_burst[1:0]         ), //i
    .io_inputs_1_payload_write (inputsCmd_1_payload_write              ), //i
    .io_inputs_2_valid         (inputsCmd_2_valid                      ), //i
    .io_inputs_2_ready         (cmdArbiter_io_inputs_2_ready           ), //o
    .io_inputs_2_payload_addr  (inputsCmd_2_payload_addr[15:0]         ), //i
    .io_inputs_2_payload_id    (inputsCmd_2_payload_id[4:0]            ), //i
    .io_inputs_2_payload_len   (inputsCmd_2_payload_len[7:0]           ), //i
    .io_inputs_2_payload_size  (inputsCmd_2_payload_size[2:0]          ), //i
    .io_inputs_2_payload_burst (inputsCmd_2_payload_burst[1:0]         ), //i
    .io_inputs_2_payload_write (inputsCmd_2_payload_write              ), //i
    .io_inputs_3_valid         (inputsCmd_3_valid                      ), //i
    .io_inputs_3_ready         (cmdArbiter_io_inputs_3_ready           ), //o
    .io_inputs_3_payload_addr  (inputsCmd_3_payload_addr[15:0]         ), //i
    .io_inputs_3_payload_id    (inputsCmd_3_payload_id[4:0]            ), //i
    .io_inputs_3_payload_len   (inputsCmd_3_payload_len[7:0]           ), //i
    .io_inputs_3_payload_size  (inputsCmd_3_payload_size[2:0]          ), //i
    .io_inputs_3_payload_burst (inputsCmd_3_payload_burst[1:0]         ), //i
    .io_inputs_3_payload_write (inputsCmd_3_payload_write              ), //i
    .io_output_valid           (cmdArbiter_io_output_valid             ), //o
    .io_output_ready           (cmdArbiter_io_output_ready             ), //i
    .io_output_payload_addr    (cmdArbiter_io_output_payload_addr[15:0]), //o
    .io_output_payload_id      (cmdArbiter_io_output_payload_id[4:0]   ), //o
    .io_output_payload_len     (cmdArbiter_io_output_payload_len[7:0]  ), //o
    .io_output_payload_size    (cmdArbiter_io_output_payload_size[2:0] ), //o
    .io_output_payload_burst   (cmdArbiter_io_output_payload_burst[1:0]), //o
    .io_output_payload_write   (cmdArbiter_io_output_payload_write     ), //o
    .io_chosen                 (cmdArbiter_io_chosen[1:0]              ), //o
    .io_chosenOH               (cmdArbiter_io_chosenOH[3:0]            ), //o
    .clk                       (clk                                    ), //i
    .reset                     (reset                                  )  //i
  );
  StreamFifoLowLatency cmdRouteFork_thrown_translated_fifo (
    .io_push_valid   (cmdRouteFork_thrown_translated_valid                    ), //i
    .io_push_ready   (cmdRouteFork_thrown_translated_fifo_io_push_ready       ), //o
    .io_push_payload (cmdRouteFork_thrown_translated_payload                  ), //i
    .io_pop_valid    (cmdRouteFork_thrown_translated_fifo_io_pop_valid        ), //o
    .io_pop_ready    (cmdRouteFork_thrown_translated_fifo_io_pop_ready        ), //i
    .io_pop_payload  (cmdRouteFork_thrown_translated_fifo_io_pop_payload      ), //o
    .io_flush        (1'b0                                                    ), //i
    .io_occupancy    (cmdRouteFork_thrown_translated_fifo_io_occupancy[2:0]   ), //o
    .io_availability (cmdRouteFork_thrown_translated_fifo_io_availability[2:0]), //o
    .clk             (clk                                                     ), //i
    .reset           (reset                                                   )  //i
  );
  always @(*) begin
    case(cmdRouteFork_thrown_translated_fifo_io_pop_payload)
      1'b0 : begin
        _zz_writeLogic_routeDataInput_valid = io_writeInputs_0_w_valid;
        _zz_writeLogic_routeDataInput_ready = io_writeInputs_0_w_ready;
        _zz_writeLogic_routeDataInput_payload_data = io_writeInputs_0_w_payload_data;
        _zz_writeLogic_routeDataInput_payload_strb = io_writeInputs_0_w_payload_strb;
        _zz_writeLogic_routeDataInput_payload_last = io_writeInputs_0_w_payload_last;
      end
      default : begin
        _zz_writeLogic_routeDataInput_valid = io_writeInputs_1_w_valid;
        _zz_writeLogic_routeDataInput_ready = io_writeInputs_1_w_ready;
        _zz_writeLogic_routeDataInput_payload_data = io_writeInputs_1_w_payload_data;
        _zz_writeLogic_routeDataInput_payload_strb = io_writeInputs_1_w_payload_strb;
        _zz_writeLogic_routeDataInput_payload_last = io_writeInputs_1_w_payload_last;
      end
    endcase
  end

  always @(*) begin
    case(writeLogic_writeRspIndex)
      1'b0 : _zz_io_output_b_ready = io_writeInputs_0_b_ready;
      default : _zz_io_output_b_ready = io_writeInputs_1_b_ready;
    endcase
  end

  always @(*) begin
    case(readRspIndex)
      1'b0 : _zz_io_output_r_ready = io_readInputs_0_r_ready;
      default : _zz_io_output_r_ready = io_readInputs_1_r_ready;
    endcase
  end

  assign inputsCmd_0_valid = io_readInputs_0_ar_valid;
  assign io_readInputs_0_ar_ready = inputsCmd_0_ready;
  assign inputsCmd_0_payload_addr = io_readInputs_0_ar_payload_addr;
  assign inputsCmd_0_payload_id = io_readInputs_0_ar_payload_id;
  assign inputsCmd_0_payload_len = io_readInputs_0_ar_payload_len;
  assign inputsCmd_0_payload_size = io_readInputs_0_ar_payload_size;
  assign inputsCmd_0_payload_burst = io_readInputs_0_ar_payload_burst;
  assign inputsCmd_0_payload_write = 1'b0;
  assign inputsCmd_1_valid = io_readInputs_1_ar_valid;
  assign io_readInputs_1_ar_ready = inputsCmd_1_ready;
  assign inputsCmd_1_payload_addr = io_readInputs_1_ar_payload_addr;
  assign inputsCmd_1_payload_id = io_readInputs_1_ar_payload_id;
  assign inputsCmd_1_payload_len = io_readInputs_1_ar_payload_len;
  assign inputsCmd_1_payload_size = io_readInputs_1_ar_payload_size;
  assign inputsCmd_1_payload_burst = io_readInputs_1_ar_payload_burst;
  assign inputsCmd_1_payload_write = 1'b0;
  assign inputsCmd_2_valid = io_writeInputs_0_aw_valid;
  assign io_writeInputs_0_aw_ready = inputsCmd_2_ready;
  assign inputsCmd_2_payload_addr = io_writeInputs_0_aw_payload_addr;
  assign inputsCmd_2_payload_id = io_writeInputs_0_aw_payload_id;
  assign inputsCmd_2_payload_len = io_writeInputs_0_aw_payload_len;
  assign inputsCmd_2_payload_size = io_writeInputs_0_aw_payload_size;
  assign inputsCmd_2_payload_burst = io_writeInputs_0_aw_payload_burst;
  assign inputsCmd_2_payload_write = 1'b1;
  assign inputsCmd_3_valid = io_writeInputs_1_aw_valid;
  assign io_writeInputs_1_aw_ready = inputsCmd_3_ready;
  assign inputsCmd_3_payload_addr = io_writeInputs_1_aw_payload_addr;
  assign inputsCmd_3_payload_id = io_writeInputs_1_aw_payload_id;
  assign inputsCmd_3_payload_len = io_writeInputs_1_aw_payload_len;
  assign inputsCmd_3_payload_size = io_writeInputs_1_aw_payload_size;
  assign inputsCmd_3_payload_burst = io_writeInputs_1_aw_payload_burst;
  assign inputsCmd_3_payload_write = 1'b1;
  assign inputsCmd_0_ready = cmdArbiter_io_inputs_0_ready;
  assign inputsCmd_1_ready = cmdArbiter_io_inputs_1_ready;
  assign inputsCmd_2_ready = cmdArbiter_io_inputs_2_ready;
  assign inputsCmd_3_ready = cmdArbiter_io_inputs_3_ready;
  always @(*) begin
    cmdArbiter_io_output_ready = 1'b1;
    if(when_Stream_l1063) begin
      cmdArbiter_io_output_ready = 1'b0;
    end
    if(when_Stream_l1063_1) begin
      cmdArbiter_io_output_ready = 1'b0;
    end
  end

  assign when_Stream_l1063 = ((! cmdOutputFork_ready) && ram_io_axi_arbiter_cmdArbiter_io_output_fork2_logic_linkEnable_0);
  assign when_Stream_l1063_1 = ((! cmdRouteFork_ready) && ram_io_axi_arbiter_cmdArbiter_io_output_fork2_logic_linkEnable_1);
  assign cmdOutputFork_valid = (cmdArbiter_io_output_valid && ram_io_axi_arbiter_cmdArbiter_io_output_fork2_logic_linkEnable_0);
  assign cmdOutputFork_payload_addr = cmdArbiter_io_output_payload_addr;
  assign cmdOutputFork_payload_id = cmdArbiter_io_output_payload_id;
  assign cmdOutputFork_payload_len = cmdArbiter_io_output_payload_len;
  assign cmdOutputFork_payload_size = cmdArbiter_io_output_payload_size;
  assign cmdOutputFork_payload_burst = cmdArbiter_io_output_payload_burst;
  assign cmdOutputFork_payload_write = cmdArbiter_io_output_payload_write;
  assign cmdOutputFork_fire = (cmdOutputFork_valid && cmdOutputFork_ready);
  assign cmdRouteFork_valid = (cmdArbiter_io_output_valid && ram_io_axi_arbiter_cmdArbiter_io_output_fork2_logic_linkEnable_1);
  assign cmdRouteFork_payload_addr = cmdArbiter_io_output_payload_addr;
  assign cmdRouteFork_payload_id = cmdArbiter_io_output_payload_id;
  assign cmdRouteFork_payload_len = cmdArbiter_io_output_payload_len;
  assign cmdRouteFork_payload_size = cmdArbiter_io_output_payload_size;
  assign cmdRouteFork_payload_burst = cmdArbiter_io_output_payload_burst;
  assign cmdRouteFork_payload_write = cmdArbiter_io_output_payload_write;
  assign cmdRouteFork_fire = (cmdRouteFork_valid && cmdRouteFork_ready);
  assign io_output_arw_valid = cmdOutputFork_valid;
  assign cmdOutputFork_ready = io_output_arw_ready;
  assign io_output_arw_payload_addr = cmdOutputFork_payload_addr;
  assign io_output_arw_payload_len = cmdOutputFork_payload_len;
  assign io_output_arw_payload_size = cmdOutputFork_payload_size;
  assign io_output_arw_payload_burst = cmdOutputFork_payload_burst;
  assign io_output_arw_payload_write = cmdOutputFork_payload_write;
  assign _zz_io_output_arw_payload_id = _zz__zz_io_output_arw_payload_id[1];
  assign _zz_io_output_arw_payload_id_1 = _zz__zz_io_output_arw_payload_id_1[1];
  assign io_output_arw_payload_id = (cmdOutputFork_payload_write ? {_zz_io_output_arw_payload_id,cmdOutputFork_payload_id} : {_zz_io_output_arw_payload_id_1,cmdOutputFork_payload_id});
  assign when_Stream_l445 = (! cmdRouteFork_payload_write);
  always @(*) begin
    cmdRouteFork_thrown_valid = cmdRouteFork_valid;
    if(when_Stream_l445) begin
      cmdRouteFork_thrown_valid = 1'b0;
    end
  end

  always @(*) begin
    cmdRouteFork_ready = cmdRouteFork_thrown_ready;
    if(when_Stream_l445) begin
      cmdRouteFork_ready = 1'b1;
    end
  end

  assign cmdRouteFork_thrown_payload_addr = cmdRouteFork_payload_addr;
  assign cmdRouteFork_thrown_payload_id = cmdRouteFork_payload_id;
  assign cmdRouteFork_thrown_payload_len = cmdRouteFork_payload_len;
  assign cmdRouteFork_thrown_payload_size = cmdRouteFork_payload_size;
  assign cmdRouteFork_thrown_payload_burst = cmdRouteFork_payload_burst;
  assign cmdRouteFork_thrown_payload_write = cmdRouteFork_payload_write;
  assign _zz_cmdRouteFork_thrown_translated_payload = _zz__zz_cmdRouteFork_thrown_translated_payload[1];
  assign cmdRouteFork_thrown_translated_valid = cmdRouteFork_thrown_valid;
  assign cmdRouteFork_thrown_ready = cmdRouteFork_thrown_translated_ready;
  assign cmdRouteFork_thrown_translated_payload = _zz_cmdRouteFork_thrown_translated_payload;
  assign cmdRouteFork_thrown_translated_ready = cmdRouteFork_thrown_translated_fifo_io_push_ready;
  assign writeLogic_routeDataInput_valid = _zz_writeLogic_routeDataInput_valid;
  assign writeLogic_routeDataInput_ready = _zz_writeLogic_routeDataInput_ready;
  assign writeLogic_routeDataInput_payload_data = _zz_writeLogic_routeDataInput_payload_data;
  assign writeLogic_routeDataInput_payload_strb = _zz_writeLogic_routeDataInput_payload_strb;
  assign writeLogic_routeDataInput_payload_last = _zz_writeLogic_routeDataInput_payload_last;
  assign io_output_w_valid = (cmdRouteFork_thrown_translated_fifo_io_pop_valid && writeLogic_routeDataInput_valid);
  assign io_output_w_payload_data = writeLogic_routeDataInput_payload_data;
  assign io_output_w_payload_strb = writeLogic_routeDataInput_payload_strb;
  assign io_output_w_payload_last = writeLogic_routeDataInput_payload_last;
  assign io_writeInputs_0_w_ready = ((cmdRouteFork_thrown_translated_fifo_io_pop_valid && io_output_w_ready) && (cmdRouteFork_thrown_translated_fifo_io_pop_payload == 1'b0));
  assign io_writeInputs_1_w_ready = ((cmdRouteFork_thrown_translated_fifo_io_pop_valid && io_output_w_ready) && (cmdRouteFork_thrown_translated_fifo_io_pop_payload == 1'b1));
  assign io_output_w_fire = (io_output_w_valid && io_output_w_ready);
  assign cmdRouteFork_thrown_translated_fifo_io_pop_ready = (io_output_w_fire && io_output_w_payload_last);
  assign writeLogic_writeRspIndex = io_output_b_payload_id[5 : 5];
  assign writeLogic_writeRspSels_0 = (writeLogic_writeRspIndex == 1'b0);
  assign writeLogic_writeRspSels_1 = (writeLogic_writeRspIndex == 1'b1);
  assign io_writeInputs_0_b_valid = (io_output_b_valid && writeLogic_writeRspSels_0);
  assign io_writeInputs_0_b_payload_resp = io_output_b_payload_resp;
  assign io_writeInputs_0_b_payload_id = io_output_b_payload_id[4:0];
  assign io_writeInputs_1_b_valid = (io_output_b_valid && writeLogic_writeRspSels_1);
  assign io_writeInputs_1_b_payload_resp = io_output_b_payload_resp;
  assign io_writeInputs_1_b_payload_id = io_output_b_payload_id[4:0];
  assign io_output_b_ready = _zz_io_output_b_ready;
  assign readRspIndex = io_output_r_payload_id[5 : 5];
  assign readRspSels_0 = (readRspIndex == 1'b0);
  assign readRspSels_1 = (readRspIndex == 1'b1);
  assign io_readInputs_0_r_valid = (io_output_r_valid && readRspSels_0);
  assign io_readInputs_0_r_payload_data = io_output_r_payload_data;
  assign io_readInputs_0_r_payload_resp = io_output_r_payload_resp;
  assign io_readInputs_0_r_payload_last = io_output_r_payload_last;
  assign io_readInputs_0_r_payload_id = io_output_r_payload_id[4:0];
  assign io_readInputs_1_r_valid = (io_output_r_valid && readRspSels_1);
  assign io_readInputs_1_r_payload_data = io_output_r_payload_data;
  assign io_readInputs_1_r_payload_resp = io_output_r_payload_resp;
  assign io_readInputs_1_r_payload_last = io_output_r_payload_last;
  assign io_readInputs_1_r_payload_id = io_output_r_payload_id[4:0];
  assign io_output_r_ready = _zz_io_output_r_ready;
  always @(posedge clk) begin
    if(reset) begin
      ram_io_axi_arbiter_cmdArbiter_io_output_fork2_logic_linkEnable_0 <= 1'b1;
      ram_io_axi_arbiter_cmdArbiter_io_output_fork2_logic_linkEnable_1 <= 1'b1;
    end else begin
      if(cmdOutputFork_fire) begin
        ram_io_axi_arbiter_cmdArbiter_io_output_fork2_logic_linkEnable_0 <= 1'b0;
      end
      if(cmdRouteFork_fire) begin
        ram_io_axi_arbiter_cmdArbiter_io_output_fork2_logic_linkEnable_1 <= 1'b0;
      end
      if(cmdArbiter_io_output_ready) begin
        ram_io_axi_arbiter_cmdArbiter_io_output_fork2_logic_linkEnable_0 <= 1'b1;
        ram_io_axi_arbiter_cmdArbiter_io_output_fork2_logic_linkEnable_1 <= 1'b1;
      end
    end
  end


endmodule

//Axi4WriteOnlyDecoder_1 replaced by Axi4WriteOnlyDecoder

//Axi4ReadOnlyDecoder_1 replaced by Axi4ReadOnlyDecoder

module Axi4WriteOnlyDecoder (
  input  wire          io_input_aw_valid,
  output wire          io_input_aw_ready,
  input  wire [31:0]   io_input_aw_payload_addr,
  input  wire [3:0]    io_input_aw_payload_id,
  input  wire [7:0]    io_input_aw_payload_len,
  input  wire [2:0]    io_input_aw_payload_size,
  input  wire [1:0]    io_input_aw_payload_burst,
  input  wire          io_input_w_valid,
  output wire          io_input_w_ready,
  input  wire [31:0]   io_input_w_payload_data,
  input  wire [3:0]    io_input_w_payload_strb,
  input  wire          io_input_w_payload_last,
  output wire          io_input_b_valid,
  input  wire          io_input_b_ready,
  output reg  [3:0]    io_input_b_payload_id,
  output reg  [1:0]    io_input_b_payload_resp,
  output wire          io_outputs_0_aw_valid,
  input  wire          io_outputs_0_aw_ready,
  output wire [31:0]   io_outputs_0_aw_payload_addr,
  output wire [3:0]    io_outputs_0_aw_payload_id,
  output wire [7:0]    io_outputs_0_aw_payload_len,
  output wire [2:0]    io_outputs_0_aw_payload_size,
  output wire [1:0]    io_outputs_0_aw_payload_burst,
  output wire          io_outputs_0_w_valid,
  input  wire          io_outputs_0_w_ready,
  output wire [31:0]   io_outputs_0_w_payload_data,
  output wire [3:0]    io_outputs_0_w_payload_strb,
  output wire          io_outputs_0_w_payload_last,
  input  wire          io_outputs_0_b_valid,
  output wire          io_outputs_0_b_ready,
  input  wire [3:0]    io_outputs_0_b_payload_id,
  input  wire [1:0]    io_outputs_0_b_payload_resp,
  input  wire          clk,
  input  wire          reset
);

  wire                errorSlave_io_axi_aw_valid;
  wire                errorSlave_io_axi_w_valid;
  wire                errorSlave_io_axi_aw_ready;
  wire                errorSlave_io_axi_w_ready;
  wire                errorSlave_io_axi_b_valid;
  wire       [3:0]    errorSlave_io_axi_b_payload_id;
  wire       [1:0]    errorSlave_io_axi_b_payload_resp;
  wire                cmdAllowedStart;
  wire                io_input_aw_fire;
  wire                io_input_b_fire;
  reg                 pendingCmdCounter_incrementIt;
  reg                 pendingCmdCounter_decrementIt;
  wire       [2:0]    pendingCmdCounter_valueNext;
  reg        [2:0]    pendingCmdCounter_value;
  wire                pendingCmdCounter_mayOverflow;
  wire                pendingCmdCounter_willOverflowIfInc;
  wire                pendingCmdCounter_willOverflow;
  reg        [2:0]    pendingCmdCounter_finalIncrement;
  wire                when_Utils_l735;
  wire                when_Utils_l737;
  wire                io_input_w_fire;
  wire                when_Utils_l709;
  reg                 pendingDataCounter_incrementIt;
  reg                 pendingDataCounter_decrementIt;
  wire       [2:0]    pendingDataCounter_valueNext;
  reg        [2:0]    pendingDataCounter_value;
  wire                pendingDataCounter_mayOverflow;
  wire                pendingDataCounter_willOverflowIfInc;
  wire                pendingDataCounter_willOverflow;
  reg        [2:0]    pendingDataCounter_finalIncrement;
  wire                when_Utils_l735_1;
  wire                when_Utils_l737_1;
  wire       [0:0]    decodedCmdSels;
  wire                decodedCmdError;
  reg        [0:0]    pendingSels;
  reg                 pendingError;
  wire                allowCmd;
  wire                allowData;
  reg                 _zz_cmdAllowedStart;

  Axi4WriteOnlyErrorSlave_1 errorSlave (
    .io_axi_aw_valid         (errorSlave_io_axi_aw_valid           ), //i
    .io_axi_aw_ready         (errorSlave_io_axi_aw_ready           ), //o
    .io_axi_aw_payload_addr  (io_input_aw_payload_addr[31:0]       ), //i
    .io_axi_aw_payload_id    (io_input_aw_payload_id[3:0]          ), //i
    .io_axi_aw_payload_len   (io_input_aw_payload_len[7:0]         ), //i
    .io_axi_aw_payload_size  (io_input_aw_payload_size[2:0]        ), //i
    .io_axi_aw_payload_burst (io_input_aw_payload_burst[1:0]       ), //i
    .io_axi_w_valid          (errorSlave_io_axi_w_valid            ), //i
    .io_axi_w_ready          (errorSlave_io_axi_w_ready            ), //o
    .io_axi_w_payload_data   (io_input_w_payload_data[31:0]        ), //i
    .io_axi_w_payload_strb   (io_input_w_payload_strb[3:0]         ), //i
    .io_axi_w_payload_last   (io_input_w_payload_last              ), //i
    .io_axi_b_valid          (errorSlave_io_axi_b_valid            ), //o
    .io_axi_b_ready          (io_input_b_ready                     ), //i
    .io_axi_b_payload_id     (errorSlave_io_axi_b_payload_id[3:0]  ), //o
    .io_axi_b_payload_resp   (errorSlave_io_axi_b_payload_resp[1:0]), //o
    .clk                     (clk                                  ), //i
    .reset                   (reset                                )  //i
  );
  assign io_input_aw_fire = (io_input_aw_valid && io_input_aw_ready);
  assign io_input_b_fire = (io_input_b_valid && io_input_b_ready);
  always @(*) begin
    pendingCmdCounter_incrementIt = 1'b0;
    if(io_input_aw_fire) begin
      pendingCmdCounter_incrementIt = 1'b1;
    end
  end

  always @(*) begin
    pendingCmdCounter_decrementIt = 1'b0;
    if(io_input_b_fire) begin
      pendingCmdCounter_decrementIt = 1'b1;
    end
  end

  assign pendingCmdCounter_mayOverflow = (pendingCmdCounter_value == 3'b111);
  assign pendingCmdCounter_willOverflowIfInc = (pendingCmdCounter_mayOverflow && (! pendingCmdCounter_decrementIt));
  assign pendingCmdCounter_willOverflow = (pendingCmdCounter_willOverflowIfInc && pendingCmdCounter_incrementIt);
  assign when_Utils_l735 = (pendingCmdCounter_incrementIt && (! pendingCmdCounter_decrementIt));
  always @(*) begin
    if(when_Utils_l735) begin
      pendingCmdCounter_finalIncrement = 3'b001;
    end else begin
      if(when_Utils_l737) begin
        pendingCmdCounter_finalIncrement = 3'b111;
      end else begin
        pendingCmdCounter_finalIncrement = 3'b000;
      end
    end
  end

  assign when_Utils_l737 = ((! pendingCmdCounter_incrementIt) && pendingCmdCounter_decrementIt);
  assign pendingCmdCounter_valueNext = (pendingCmdCounter_value + pendingCmdCounter_finalIncrement);
  assign io_input_w_fire = (io_input_w_valid && io_input_w_ready);
  assign when_Utils_l709 = (io_input_w_fire && io_input_w_payload_last);
  always @(*) begin
    pendingDataCounter_incrementIt = 1'b0;
    if(cmdAllowedStart) begin
      pendingDataCounter_incrementIt = 1'b1;
    end
  end

  always @(*) begin
    pendingDataCounter_decrementIt = 1'b0;
    if(when_Utils_l709) begin
      pendingDataCounter_decrementIt = 1'b1;
    end
  end

  assign pendingDataCounter_mayOverflow = (pendingDataCounter_value == 3'b111);
  assign pendingDataCounter_willOverflowIfInc = (pendingDataCounter_mayOverflow && (! pendingDataCounter_decrementIt));
  assign pendingDataCounter_willOverflow = (pendingDataCounter_willOverflowIfInc && pendingDataCounter_incrementIt);
  assign when_Utils_l735_1 = (pendingDataCounter_incrementIt && (! pendingDataCounter_decrementIt));
  always @(*) begin
    if(when_Utils_l735_1) begin
      pendingDataCounter_finalIncrement = 3'b001;
    end else begin
      if(when_Utils_l737_1) begin
        pendingDataCounter_finalIncrement = 3'b111;
      end else begin
        pendingDataCounter_finalIncrement = 3'b000;
      end
    end
  end

  assign when_Utils_l737_1 = ((! pendingDataCounter_incrementIt) && pendingDataCounter_decrementIt);
  assign pendingDataCounter_valueNext = (pendingDataCounter_value + pendingDataCounter_finalIncrement);
  assign decodedCmdSels = (((io_input_aw_payload_addr & (~ 32'h0000ffff)) == 32'h0) && io_input_aw_valid);
  assign decodedCmdError = (decodedCmdSels == 1'b0);
  assign allowCmd = ((pendingCmdCounter_value == 3'b000) || ((pendingCmdCounter_value != 3'b111) && (pendingSels == decodedCmdSels)));
  assign allowData = (pendingDataCounter_value != 3'b000);
  assign cmdAllowedStart = ((io_input_aw_valid && allowCmd) && _zz_cmdAllowedStart);
  assign io_input_aw_ready = (((|(decodedCmdSels & io_outputs_0_aw_ready)) || (decodedCmdError && errorSlave_io_axi_aw_ready)) && allowCmd);
  assign errorSlave_io_axi_aw_valid = ((io_input_aw_valid && decodedCmdError) && allowCmd);
  assign io_outputs_0_aw_valid = ((io_input_aw_valid && decodedCmdSels[0]) && allowCmd);
  assign io_outputs_0_aw_payload_addr = io_input_aw_payload_addr;
  assign io_outputs_0_aw_payload_id = io_input_aw_payload_id;
  assign io_outputs_0_aw_payload_len = io_input_aw_payload_len;
  assign io_outputs_0_aw_payload_size = io_input_aw_payload_size;
  assign io_outputs_0_aw_payload_burst = io_input_aw_payload_burst;
  assign io_input_w_ready = (((|(pendingSels & io_outputs_0_w_ready)) || (pendingError && errorSlave_io_axi_w_ready)) && allowData);
  assign errorSlave_io_axi_w_valid = ((io_input_w_valid && pendingError) && allowData);
  assign io_outputs_0_w_valid = ((io_input_w_valid && pendingSels[0]) && allowData);
  assign io_outputs_0_w_payload_data = io_input_w_payload_data;
  assign io_outputs_0_w_payload_strb = io_input_w_payload_strb;
  assign io_outputs_0_w_payload_last = io_input_w_payload_last;
  assign io_input_b_valid = ((|io_outputs_0_b_valid) || errorSlave_io_axi_b_valid);
  always @(*) begin
    io_input_b_payload_id = io_outputs_0_b_payload_id;
    if(pendingError) begin
      io_input_b_payload_id = errorSlave_io_axi_b_payload_id;
    end
  end

  always @(*) begin
    io_input_b_payload_resp = io_outputs_0_b_payload_resp;
    if(pendingError) begin
      io_input_b_payload_resp = errorSlave_io_axi_b_payload_resp;
    end
  end

  assign io_outputs_0_b_ready = io_input_b_ready;
  always @(posedge clk) begin
    if(reset) begin
      pendingCmdCounter_value <= 3'b000;
      pendingDataCounter_value <= 3'b000;
      pendingSels <= 1'b0;
      pendingError <= 1'b0;
      _zz_cmdAllowedStart <= 1'b1;
    end else begin
      pendingCmdCounter_value <= pendingCmdCounter_valueNext;
      pendingDataCounter_value <= pendingDataCounter_valueNext;
      if(cmdAllowedStart) begin
        pendingSels <= decodedCmdSels;
      end
      if(cmdAllowedStart) begin
        pendingError <= decodedCmdError;
      end
      if(cmdAllowedStart) begin
        _zz_cmdAllowedStart <= 1'b0;
      end
      if(io_input_aw_ready) begin
        _zz_cmdAllowedStart <= 1'b1;
      end
    end
  end


endmodule

module Axi4ReadOnlyDecoder (
  input  wire          io_input_ar_valid,
  output wire          io_input_ar_ready,
  input  wire [31:0]   io_input_ar_payload_addr,
  input  wire [3:0]    io_input_ar_payload_id,
  input  wire [7:0]    io_input_ar_payload_len,
  input  wire [2:0]    io_input_ar_payload_size,
  input  wire [1:0]    io_input_ar_payload_burst,
  output reg           io_input_r_valid,
  input  wire          io_input_r_ready,
  output wire [31:0]   io_input_r_payload_data,
  output reg  [3:0]    io_input_r_payload_id,
  output reg  [1:0]    io_input_r_payload_resp,
  output reg           io_input_r_payload_last,
  output wire          io_outputs_0_ar_valid,
  input  wire          io_outputs_0_ar_ready,
  output wire [31:0]   io_outputs_0_ar_payload_addr,
  output wire [3:0]    io_outputs_0_ar_payload_id,
  output wire [7:0]    io_outputs_0_ar_payload_len,
  output wire [2:0]    io_outputs_0_ar_payload_size,
  output wire [1:0]    io_outputs_0_ar_payload_burst,
  input  wire          io_outputs_0_r_valid,
  output wire          io_outputs_0_r_ready,
  input  wire [31:0]   io_outputs_0_r_payload_data,
  input  wire [3:0]    io_outputs_0_r_payload_id,
  input  wire [1:0]    io_outputs_0_r_payload_resp,
  input  wire          io_outputs_0_r_payload_last,
  input  wire          clk,
  input  wire          reset
);

  wire                errorSlave_io_axi_ar_valid;
  wire                errorSlave_io_axi_ar_ready;
  wire                errorSlave_io_axi_r_valid;
  wire       [31:0]   errorSlave_io_axi_r_payload_data;
  wire       [3:0]    errorSlave_io_axi_r_payload_id;
  wire       [1:0]    errorSlave_io_axi_r_payload_resp;
  wire                errorSlave_io_axi_r_payload_last;
  wire                io_input_ar_fire;
  wire                io_input_r_fire;
  wire                when_Utils_l709;
  reg                 pendingCmdCounter_incrementIt;
  reg                 pendingCmdCounter_decrementIt;
  wire       [2:0]    pendingCmdCounter_valueNext;
  reg        [2:0]    pendingCmdCounter_value;
  wire                pendingCmdCounter_mayOverflow;
  wire                pendingCmdCounter_willOverflowIfInc;
  wire                pendingCmdCounter_willOverflow;
  reg        [2:0]    pendingCmdCounter_finalIncrement;
  wire                when_Utils_l735;
  wire                when_Utils_l737;
  wire       [0:0]    decodedCmdSels;
  wire                decodedCmdError;
  reg        [0:0]    pendingSels;
  reg                 pendingError;
  wire                allowCmd;

  Axi4ReadOnlyErrorSlave_1 errorSlave (
    .io_axi_ar_valid         (errorSlave_io_axi_ar_valid            ), //i
    .io_axi_ar_ready         (errorSlave_io_axi_ar_ready            ), //o
    .io_axi_ar_payload_addr  (io_input_ar_payload_addr[31:0]        ), //i
    .io_axi_ar_payload_id    (io_input_ar_payload_id[3:0]           ), //i
    .io_axi_ar_payload_len   (io_input_ar_payload_len[7:0]          ), //i
    .io_axi_ar_payload_size  (io_input_ar_payload_size[2:0]         ), //i
    .io_axi_ar_payload_burst (io_input_ar_payload_burst[1:0]        ), //i
    .io_axi_r_valid          (errorSlave_io_axi_r_valid             ), //o
    .io_axi_r_ready          (io_input_r_ready                      ), //i
    .io_axi_r_payload_data   (errorSlave_io_axi_r_payload_data[31:0]), //o
    .io_axi_r_payload_id     (errorSlave_io_axi_r_payload_id[3:0]   ), //o
    .io_axi_r_payload_resp   (errorSlave_io_axi_r_payload_resp[1:0] ), //o
    .io_axi_r_payload_last   (errorSlave_io_axi_r_payload_last      ), //o
    .clk                     (clk                                   ), //i
    .reset                   (reset                                 )  //i
  );
  assign io_input_ar_fire = (io_input_ar_valid && io_input_ar_ready);
  assign io_input_r_fire = (io_input_r_valid && io_input_r_ready);
  assign when_Utils_l709 = (io_input_r_fire && io_input_r_payload_last);
  always @(*) begin
    pendingCmdCounter_incrementIt = 1'b0;
    if(io_input_ar_fire) begin
      pendingCmdCounter_incrementIt = 1'b1;
    end
  end

  always @(*) begin
    pendingCmdCounter_decrementIt = 1'b0;
    if(when_Utils_l709) begin
      pendingCmdCounter_decrementIt = 1'b1;
    end
  end

  assign pendingCmdCounter_mayOverflow = (pendingCmdCounter_value == 3'b111);
  assign pendingCmdCounter_willOverflowIfInc = (pendingCmdCounter_mayOverflow && (! pendingCmdCounter_decrementIt));
  assign pendingCmdCounter_willOverflow = (pendingCmdCounter_willOverflowIfInc && pendingCmdCounter_incrementIt);
  assign when_Utils_l735 = (pendingCmdCounter_incrementIt && (! pendingCmdCounter_decrementIt));
  always @(*) begin
    if(when_Utils_l735) begin
      pendingCmdCounter_finalIncrement = 3'b001;
    end else begin
      if(when_Utils_l737) begin
        pendingCmdCounter_finalIncrement = 3'b111;
      end else begin
        pendingCmdCounter_finalIncrement = 3'b000;
      end
    end
  end

  assign when_Utils_l737 = ((! pendingCmdCounter_incrementIt) && pendingCmdCounter_decrementIt);
  assign pendingCmdCounter_valueNext = (pendingCmdCounter_value + pendingCmdCounter_finalIncrement);
  assign decodedCmdSels = (((io_input_ar_payload_addr & (~ 32'h0000ffff)) == 32'h0) && io_input_ar_valid);
  assign decodedCmdError = (decodedCmdSels == 1'b0);
  assign allowCmd = ((pendingCmdCounter_value == 3'b000) || ((pendingCmdCounter_value != 3'b111) && (pendingSels == decodedCmdSels)));
  assign io_input_ar_ready = (((|(decodedCmdSels & io_outputs_0_ar_ready)) || (decodedCmdError && errorSlave_io_axi_ar_ready)) && allowCmd);
  assign errorSlave_io_axi_ar_valid = ((io_input_ar_valid && decodedCmdError) && allowCmd);
  assign io_outputs_0_ar_valid = ((io_input_ar_valid && decodedCmdSels[0]) && allowCmd);
  assign io_outputs_0_ar_payload_addr = io_input_ar_payload_addr;
  assign io_outputs_0_ar_payload_id = io_input_ar_payload_id;
  assign io_outputs_0_ar_payload_len = io_input_ar_payload_len;
  assign io_outputs_0_ar_payload_size = io_input_ar_payload_size;
  assign io_outputs_0_ar_payload_burst = io_input_ar_payload_burst;
  always @(*) begin
    io_input_r_valid = (|io_outputs_0_r_valid);
    if(errorSlave_io_axi_r_valid) begin
      io_input_r_valid = 1'b1;
    end
  end

  assign io_input_r_payload_data = io_outputs_0_r_payload_data;
  always @(*) begin
    io_input_r_payload_id = io_outputs_0_r_payload_id;
    if(pendingError) begin
      io_input_r_payload_id = errorSlave_io_axi_r_payload_id;
    end
  end

  always @(*) begin
    io_input_r_payload_resp = io_outputs_0_r_payload_resp;
    if(pendingError) begin
      io_input_r_payload_resp = errorSlave_io_axi_r_payload_resp;
    end
  end

  always @(*) begin
    io_input_r_payload_last = io_outputs_0_r_payload_last;
    if(pendingError) begin
      io_input_r_payload_last = errorSlave_io_axi_r_payload_last;
    end
  end

  assign io_outputs_0_r_ready = io_input_r_ready;
  always @(posedge clk) begin
    if(reset) begin
      pendingCmdCounter_value <= 3'b000;
      pendingSels <= 1'b0;
      pendingError <= 1'b0;
    end else begin
      pendingCmdCounter_value <= pendingCmdCounter_valueNext;
      if(io_input_ar_ready) begin
        pendingSels <= decodedCmdSels;
      end
      if(io_input_ar_ready) begin
        pendingError <= decodedCmdError;
      end
    end
  end


endmodule

module Axi4SharedOnChipRam (
  input  wire          io_axi_arw_valid,
  output wire          io_axi_arw_ready,
  input  wire [15:0]   io_axi_arw_payload_addr,
  input  wire [5:0]    io_axi_arw_payload_id,
  input  wire [7:0]    io_axi_arw_payload_len,
  input  wire [2:0]    io_axi_arw_payload_size,
  input  wire [1:0]    io_axi_arw_payload_burst,
  input  wire          io_axi_arw_payload_write,
  input  wire          io_axi_w_valid,
  output wire          io_axi_w_ready,
  input  wire [31:0]   io_axi_w_payload_data,
  input  wire [3:0]    io_axi_w_payload_strb,
  input  wire          io_axi_w_payload_last,
  output wire          io_axi_b_valid,
  input  wire          io_axi_b_ready,
  output wire [5:0]    io_axi_b_payload_id,
  output wire [1:0]    io_axi_b_payload_resp,
  output wire          io_axi_r_valid,
  input  wire          io_axi_r_ready,
  output wire [31:0]   io_axi_r_payload_data,
  output wire [5:0]    io_axi_r_payload_id,
  output wire [1:0]    io_axi_r_payload_resp,
  output wire          io_axi_r_payload_last,
  input  wire          clk,
  input  wire          reset
);

  reg        [31:0]   ram_spinal_port0;
  wire       [1:0]    _zz_Axi4Incr_alignMask;
  wire       [11:0]   _zz_Axi4Incr_baseIncr;
  wire       [2:0]    _zz_Axi4Incr_wrapCase_1;
  wire       [2:0]    _zz_Axi4Incr_wrapCase_2;
  reg        [11:0]   _zz_Axi4Incr_result;
  wire       [10:0]   _zz_Axi4Incr_result_1;
  wire       [0:0]    _zz_Axi4Incr_result_2;
  wire       [9:0]    _zz_Axi4Incr_result_3;
  wire       [1:0]    _zz_Axi4Incr_result_4;
  wire       [8:0]    _zz_Axi4Incr_result_5;
  wire       [2:0]    _zz_Axi4Incr_result_6;
  wire       [7:0]    _zz_Axi4Incr_result_7;
  wire       [3:0]    _zz_Axi4Incr_result_8;
  wire       [6:0]    _zz_Axi4Incr_result_9;
  wire       [4:0]    _zz_Axi4Incr_result_10;
  wire       [5:0]    _zz_Axi4Incr_result_11;
  wire       [5:0]    _zz_Axi4Incr_result_12;
  wire                io_axi_arw_s2mPipe_valid;
  reg                 io_axi_arw_s2mPipe_ready;
  wire       [15:0]   io_axi_arw_s2mPipe_payload_addr;
  wire       [5:0]    io_axi_arw_s2mPipe_payload_id;
  wire       [7:0]    io_axi_arw_s2mPipe_payload_len;
  wire       [2:0]    io_axi_arw_s2mPipe_payload_size;
  wire       [1:0]    io_axi_arw_s2mPipe_payload_burst;
  wire                io_axi_arw_s2mPipe_payload_write;
  reg                 io_axi_arw_rValidN;
  reg        [15:0]   io_axi_arw_rData_addr;
  reg        [5:0]    io_axi_arw_rData_id;
  reg        [7:0]    io_axi_arw_rData_len;
  reg        [2:0]    io_axi_arw_rData_size;
  reg        [1:0]    io_axi_arw_rData_burst;
  reg                 io_axi_arw_rData_write;
  reg                 unburstify_result_valid;
  reg                 unburstify_result_ready;
  reg                 unburstify_result_payload_last;
  reg        [15:0]   unburstify_result_payload_fragment_addr;
  reg        [5:0]    unburstify_result_payload_fragment_id;
  reg        [2:0]    unburstify_result_payload_fragment_size;
  reg        [1:0]    unburstify_result_payload_fragment_burst;
  reg                 unburstify_result_payload_fragment_write;
  wire                unburstify_doResult;
  reg                 unburstify_buffer_valid;
  reg        [7:0]    unburstify_buffer_len;
  reg        [7:0]    unburstify_buffer_beat;
  reg        [15:0]   unburstify_buffer_transaction_addr;
  reg        [5:0]    unburstify_buffer_transaction_id;
  reg        [2:0]    unburstify_buffer_transaction_size;
  reg        [1:0]    unburstify_buffer_transaction_burst;
  reg                 unburstify_buffer_transaction_write;
  wire                unburstify_buffer_last;
  wire       [1:0]    Axi4Incr_validSize;
  reg        [15:0]   Axi4Incr_result;
  wire       [3:0]    Axi4Incr_highCat;
  wire       [2:0]    Axi4Incr_sizeValue;
  wire       [11:0]   Axi4Incr_alignMask;
  wire       [11:0]   Axi4Incr_base;
  wire       [11:0]   Axi4Incr_baseIncr;
  reg        [1:0]    _zz_Axi4Incr_wrapCase;
  wire       [2:0]    Axi4Incr_wrapCase;
  wire                when_Axi4Channel_l322;
  wire                arw_valid;
  wire                arw_ready;
  wire                arw_payload_last;
  wire       [15:0]   arw_payload_fragment_addr;
  wire       [5:0]    arw_payload_fragment_id;
  wire       [2:0]    arw_payload_fragment_size;
  wire       [1:0]    arw_payload_fragment_burst;
  wire                arw_payload_fragment_write;
  reg                 unburstify_result_rValid;
  reg                 unburstify_result_rData_last;
  reg        [15:0]   unburstify_result_rData_fragment_addr;
  reg        [5:0]    unburstify_result_rData_fragment_id;
  reg        [2:0]    unburstify_result_rData_fragment_size;
  reg        [1:0]    unburstify_result_rData_fragment_burst;
  reg                 unburstify_result_rData_fragment_write;
  wire                when_Stream_l375;
  wire                _zz_arw_ready;
  wire                stage0_valid;
  reg                 stage0_ready;
  wire                stage0_payload_last;
  wire       [15:0]   stage0_payload_fragment_addr;
  wire       [5:0]    stage0_payload_fragment_id;
  wire       [2:0]    stage0_payload_fragment_size;
  wire       [1:0]    stage0_payload_fragment_burst;
  wire                stage0_payload_fragment_write;
  wire       [13:0]   _zz_io_axi_r_payload_data;
  wire                stage0_fire;
  wire       [31:0]   _zz_io_axi_r_payload_data_1;
  wire                stage1_valid;
  wire                stage1_ready;
  wire                stage1_payload_last;
  wire       [15:0]   stage1_payload_fragment_addr;
  wire       [5:0]    stage1_payload_fragment_id;
  wire       [2:0]    stage1_payload_fragment_size;
  wire       [1:0]    stage1_payload_fragment_burst;
  wire                stage1_payload_fragment_write;
  reg                 stage0_rValid;
  reg                 stage0_rData_last;
  reg        [15:0]   stage0_rData_fragment_addr;
  reg        [5:0]    stage0_rData_fragment_id;
  reg        [2:0]    stage0_rData_fragment_size;
  reg        [1:0]    stage0_rData_fragment_burst;
  reg                 stage0_rData_fragment_write;
  wire                when_Stream_l375_1;
  reg [7:0] ram_symbol0 [0:16383];
  reg [7:0] ram_symbol1 [0:16383];
  reg [7:0] ram_symbol2 [0:16383];
  reg [7:0] ram_symbol3 [0:16383];
  reg [7:0] _zz_ramsymbol_read;
  reg [7:0] _zz_ramsymbol_read_1;
  reg [7:0] _zz_ramsymbol_read_2;
  reg [7:0] _zz_ramsymbol_read_3;

  assign _zz_Axi4Incr_alignMask = {(2'b01 < Axi4Incr_validSize),(2'b00 < Axi4Incr_validSize)};
  assign _zz_Axi4Incr_baseIncr = {9'd0, Axi4Incr_sizeValue};
  assign _zz_Axi4Incr_wrapCase_1 = {1'd0, Axi4Incr_validSize};
  assign _zz_Axi4Incr_wrapCase_2 = {1'd0, _zz_Axi4Incr_wrapCase};
  assign _zz_Axi4Incr_result_1 = Axi4Incr_base[11 : 1];
  assign _zz_Axi4Incr_result_2 = Axi4Incr_baseIncr[0 : 0];
  assign _zz_Axi4Incr_result_3 = Axi4Incr_base[11 : 2];
  assign _zz_Axi4Incr_result_4 = Axi4Incr_baseIncr[1 : 0];
  assign _zz_Axi4Incr_result_5 = Axi4Incr_base[11 : 3];
  assign _zz_Axi4Incr_result_6 = Axi4Incr_baseIncr[2 : 0];
  assign _zz_Axi4Incr_result_7 = Axi4Incr_base[11 : 4];
  assign _zz_Axi4Incr_result_8 = Axi4Incr_baseIncr[3 : 0];
  assign _zz_Axi4Incr_result_9 = Axi4Incr_base[11 : 5];
  assign _zz_Axi4Incr_result_10 = Axi4Incr_baseIncr[4 : 0];
  assign _zz_Axi4Incr_result_11 = Axi4Incr_base[11 : 6];
  assign _zz_Axi4Incr_result_12 = Axi4Incr_baseIncr[5 : 0];
  always @(*) begin
    ram_spinal_port0 = {_zz_ramsymbol_read_3, _zz_ramsymbol_read_2, _zz_ramsymbol_read_1, _zz_ramsymbol_read};
  end
  always @(posedge clk) begin
    if(stage0_fire) begin
      _zz_ramsymbol_read <= ram_symbol0[_zz_io_axi_r_payload_data];
      _zz_ramsymbol_read_1 <= ram_symbol1[_zz_io_axi_r_payload_data];
      _zz_ramsymbol_read_2 <= ram_symbol2[_zz_io_axi_r_payload_data];
      _zz_ramsymbol_read_3 <= ram_symbol3[_zz_io_axi_r_payload_data];
    end
  end

  always @(posedge clk) begin
    if(io_axi_w_payload_strb[0] && stage0_fire && stage0_payload_fragment_write ) begin
      ram_symbol0[_zz_io_axi_r_payload_data] <= _zz_io_axi_r_payload_data_1[7 : 0];
    end
    if(io_axi_w_payload_strb[1] && stage0_fire && stage0_payload_fragment_write ) begin
      ram_symbol1[_zz_io_axi_r_payload_data] <= _zz_io_axi_r_payload_data_1[15 : 8];
    end
    if(io_axi_w_payload_strb[2] && stage0_fire && stage0_payload_fragment_write ) begin
      ram_symbol2[_zz_io_axi_r_payload_data] <= _zz_io_axi_r_payload_data_1[23 : 16];
    end
    if(io_axi_w_payload_strb[3] && stage0_fire && stage0_payload_fragment_write ) begin
      ram_symbol3[_zz_io_axi_r_payload_data] <= _zz_io_axi_r_payload_data_1[31 : 24];
    end
  end

  always @(*) begin
    case(Axi4Incr_wrapCase)
      3'b000 : _zz_Axi4Incr_result = {_zz_Axi4Incr_result_1,_zz_Axi4Incr_result_2};
      3'b001 : _zz_Axi4Incr_result = {_zz_Axi4Incr_result_3,_zz_Axi4Incr_result_4};
      3'b010 : _zz_Axi4Incr_result = {_zz_Axi4Incr_result_5,_zz_Axi4Incr_result_6};
      3'b011 : _zz_Axi4Incr_result = {_zz_Axi4Incr_result_7,_zz_Axi4Incr_result_8};
      3'b100 : _zz_Axi4Incr_result = {_zz_Axi4Incr_result_9,_zz_Axi4Incr_result_10};
      default : _zz_Axi4Incr_result = {_zz_Axi4Incr_result_11,_zz_Axi4Incr_result_12};
    endcase
  end

  assign io_axi_arw_ready = io_axi_arw_rValidN;
  assign io_axi_arw_s2mPipe_valid = (io_axi_arw_valid || (! io_axi_arw_rValidN));
  assign io_axi_arw_s2mPipe_payload_addr = (io_axi_arw_rValidN ? io_axi_arw_payload_addr : io_axi_arw_rData_addr);
  assign io_axi_arw_s2mPipe_payload_id = (io_axi_arw_rValidN ? io_axi_arw_payload_id : io_axi_arw_rData_id);
  assign io_axi_arw_s2mPipe_payload_len = (io_axi_arw_rValidN ? io_axi_arw_payload_len : io_axi_arw_rData_len);
  assign io_axi_arw_s2mPipe_payload_size = (io_axi_arw_rValidN ? io_axi_arw_payload_size : io_axi_arw_rData_size);
  assign io_axi_arw_s2mPipe_payload_burst = (io_axi_arw_rValidN ? io_axi_arw_payload_burst : io_axi_arw_rData_burst);
  assign io_axi_arw_s2mPipe_payload_write = (io_axi_arw_rValidN ? io_axi_arw_payload_write : io_axi_arw_rData_write);
  assign unburstify_buffer_last = (unburstify_buffer_beat == 8'h01);
  assign Axi4Incr_validSize = unburstify_buffer_transaction_size[1 : 0];
  assign Axi4Incr_highCat = unburstify_buffer_transaction_addr[15 : 12];
  assign Axi4Incr_sizeValue = {(2'b10 == Axi4Incr_validSize),{(2'b01 == Axi4Incr_validSize),(2'b00 == Axi4Incr_validSize)}};
  assign Axi4Incr_alignMask = {10'd0, _zz_Axi4Incr_alignMask};
  assign Axi4Incr_base = (unburstify_buffer_transaction_addr[11 : 0] & (~ Axi4Incr_alignMask));
  assign Axi4Incr_baseIncr = (Axi4Incr_base + _zz_Axi4Incr_baseIncr);
  always @(*) begin
    casez(unburstify_buffer_len)
      8'b????1??? : begin
        _zz_Axi4Incr_wrapCase = 2'b11;
      end
      8'b????01?? : begin
        _zz_Axi4Incr_wrapCase = 2'b10;
      end
      8'b????001? : begin
        _zz_Axi4Incr_wrapCase = 2'b01;
      end
      default : begin
        _zz_Axi4Incr_wrapCase = 2'b00;
      end
    endcase
  end

  assign Axi4Incr_wrapCase = (_zz_Axi4Incr_wrapCase_1 + _zz_Axi4Incr_wrapCase_2);
  always @(*) begin
    case(unburstify_buffer_transaction_burst)
      2'b00 : begin
        Axi4Incr_result = unburstify_buffer_transaction_addr;
      end
      2'b10 : begin
        Axi4Incr_result = {Axi4Incr_highCat,_zz_Axi4Incr_result};
      end
      default : begin
        Axi4Incr_result = {Axi4Incr_highCat,Axi4Incr_baseIncr};
      end
    endcase
  end

  always @(*) begin
    io_axi_arw_s2mPipe_ready = 1'b0;
    if(!unburstify_buffer_valid) begin
      io_axi_arw_s2mPipe_ready = unburstify_result_ready;
    end
  end

  always @(*) begin
    if(unburstify_buffer_valid) begin
      unburstify_result_valid = 1'b1;
    end else begin
      unburstify_result_valid = io_axi_arw_s2mPipe_valid;
    end
  end

  always @(*) begin
    if(unburstify_buffer_valid) begin
      unburstify_result_payload_last = unburstify_buffer_last;
    end else begin
      unburstify_result_payload_last = 1'b1;
      if(when_Axi4Channel_l322) begin
        unburstify_result_payload_last = 1'b0;
      end
    end
  end

  always @(*) begin
    if(unburstify_buffer_valid) begin
      unburstify_result_payload_fragment_id = unburstify_buffer_transaction_id;
    end else begin
      unburstify_result_payload_fragment_id = io_axi_arw_s2mPipe_payload_id;
    end
  end

  always @(*) begin
    if(unburstify_buffer_valid) begin
      unburstify_result_payload_fragment_size = unburstify_buffer_transaction_size;
    end else begin
      unburstify_result_payload_fragment_size = io_axi_arw_s2mPipe_payload_size;
    end
  end

  always @(*) begin
    if(unburstify_buffer_valid) begin
      unburstify_result_payload_fragment_burst = unburstify_buffer_transaction_burst;
    end else begin
      unburstify_result_payload_fragment_burst = io_axi_arw_s2mPipe_payload_burst;
    end
  end

  always @(*) begin
    if(unburstify_buffer_valid) begin
      unburstify_result_payload_fragment_write = unburstify_buffer_transaction_write;
    end else begin
      unburstify_result_payload_fragment_write = io_axi_arw_s2mPipe_payload_write;
    end
  end

  always @(*) begin
    if(unburstify_buffer_valid) begin
      unburstify_result_payload_fragment_addr = Axi4Incr_result;
    end else begin
      unburstify_result_payload_fragment_addr = io_axi_arw_s2mPipe_payload_addr;
    end
  end

  assign when_Axi4Channel_l322 = (io_axi_arw_s2mPipe_payload_len != 8'h0);
  always @(*) begin
    unburstify_result_ready = arw_ready;
    if(when_Stream_l375) begin
      unburstify_result_ready = 1'b1;
    end
  end

  assign when_Stream_l375 = (! arw_valid);
  assign arw_valid = unburstify_result_rValid;
  assign arw_payload_last = unburstify_result_rData_last;
  assign arw_payload_fragment_addr = unburstify_result_rData_fragment_addr;
  assign arw_payload_fragment_id = unburstify_result_rData_fragment_id;
  assign arw_payload_fragment_size = unburstify_result_rData_fragment_size;
  assign arw_payload_fragment_burst = unburstify_result_rData_fragment_burst;
  assign arw_payload_fragment_write = unburstify_result_rData_fragment_write;
  assign _zz_arw_ready = (! (arw_payload_fragment_write && (! io_axi_w_valid)));
  assign stage0_valid = (arw_valid && _zz_arw_ready);
  assign arw_ready = (stage0_ready && _zz_arw_ready);
  assign stage0_payload_last = arw_payload_last;
  assign stage0_payload_fragment_addr = arw_payload_fragment_addr;
  assign stage0_payload_fragment_id = arw_payload_fragment_id;
  assign stage0_payload_fragment_size = arw_payload_fragment_size;
  assign stage0_payload_fragment_burst = arw_payload_fragment_burst;
  assign stage0_payload_fragment_write = arw_payload_fragment_write;
  assign _zz_io_axi_r_payload_data = stage0_payload_fragment_addr[15 : 2];
  assign stage0_fire = (stage0_valid && stage0_ready);
  assign _zz_io_axi_r_payload_data_1 = io_axi_w_payload_data;
  assign io_axi_r_payload_data = ram_spinal_port0;
  assign io_axi_w_ready = ((arw_valid && arw_payload_fragment_write) && stage0_ready);
  always @(*) begin
    stage0_ready = stage1_ready;
    if(when_Stream_l375_1) begin
      stage0_ready = 1'b1;
    end
  end

  assign when_Stream_l375_1 = (! stage1_valid);
  assign stage1_valid = stage0_rValid;
  assign stage1_payload_last = stage0_rData_last;
  assign stage1_payload_fragment_addr = stage0_rData_fragment_addr;
  assign stage1_payload_fragment_id = stage0_rData_fragment_id;
  assign stage1_payload_fragment_size = stage0_rData_fragment_size;
  assign stage1_payload_fragment_burst = stage0_rData_fragment_burst;
  assign stage1_payload_fragment_write = stage0_rData_fragment_write;
  assign stage1_ready = ((io_axi_r_ready && (! stage1_payload_fragment_write)) || ((io_axi_b_ready || (! stage1_payload_last)) && stage1_payload_fragment_write));
  assign io_axi_r_valid = (stage1_valid && (! stage1_payload_fragment_write));
  assign io_axi_r_payload_id = stage1_payload_fragment_id;
  assign io_axi_r_payload_last = stage1_payload_last;
  assign io_axi_r_payload_resp = 2'b00;
  assign io_axi_b_valid = ((stage1_valid && stage1_payload_fragment_write) && stage1_payload_last);
  assign io_axi_b_payload_resp = 2'b00;
  assign io_axi_b_payload_id = stage1_payload_fragment_id;
  always @(posedge clk) begin
    if(reset) begin
      io_axi_arw_rValidN <= 1'b1;
      unburstify_buffer_valid <= 1'b0;
      unburstify_result_rValid <= 1'b0;
      stage0_rValid <= 1'b0;
    end else begin
      if(io_axi_arw_valid) begin
        io_axi_arw_rValidN <= 1'b0;
      end
      if(io_axi_arw_s2mPipe_ready) begin
        io_axi_arw_rValidN <= 1'b1;
      end
      if(unburstify_result_ready) begin
        if(unburstify_buffer_last) begin
          unburstify_buffer_valid <= 1'b0;
        end
      end
      if(!unburstify_buffer_valid) begin
        if(when_Axi4Channel_l322) begin
          if(unburstify_result_ready) begin
            unburstify_buffer_valid <= io_axi_arw_s2mPipe_valid;
          end
        end
      end
      if(unburstify_result_ready) begin
        unburstify_result_rValid <= unburstify_result_valid;
      end
      if(stage0_ready) begin
        stage0_rValid <= stage0_valid;
      end
    end
  end

  always @(posedge clk) begin
    if(io_axi_arw_ready) begin
      io_axi_arw_rData_addr <= io_axi_arw_payload_addr;
      io_axi_arw_rData_id <= io_axi_arw_payload_id;
      io_axi_arw_rData_len <= io_axi_arw_payload_len;
      io_axi_arw_rData_size <= io_axi_arw_payload_size;
      io_axi_arw_rData_burst <= io_axi_arw_payload_burst;
      io_axi_arw_rData_write <= io_axi_arw_payload_write;
    end
    if(unburstify_result_ready) begin
      unburstify_buffer_beat <= (unburstify_buffer_beat - 8'h01);
      unburstify_buffer_transaction_addr[11 : 0] <= Axi4Incr_result[11 : 0];
    end
    if(!unburstify_buffer_valid) begin
      if(when_Axi4Channel_l322) begin
        if(unburstify_result_ready) begin
          unburstify_buffer_transaction_addr <= io_axi_arw_s2mPipe_payload_addr;
          unburstify_buffer_transaction_id <= io_axi_arw_s2mPipe_payload_id;
          unburstify_buffer_transaction_size <= io_axi_arw_s2mPipe_payload_size;
          unburstify_buffer_transaction_burst <= io_axi_arw_s2mPipe_payload_burst;
          unburstify_buffer_transaction_write <= io_axi_arw_s2mPipe_payload_write;
          unburstify_buffer_beat <= io_axi_arw_s2mPipe_payload_len;
          unburstify_buffer_len <= io_axi_arw_s2mPipe_payload_len;
        end
      end
    end
    if(unburstify_result_ready) begin
      unburstify_result_rData_last <= unburstify_result_payload_last;
      unburstify_result_rData_fragment_addr <= unburstify_result_payload_fragment_addr;
      unburstify_result_rData_fragment_id <= unburstify_result_payload_fragment_id;
      unburstify_result_rData_fragment_size <= unburstify_result_payload_fragment_size;
      unburstify_result_rData_fragment_burst <= unburstify_result_payload_fragment_burst;
      unburstify_result_rData_fragment_write <= unburstify_result_payload_fragment_write;
    end
    if(stage0_ready) begin
      stage0_rData_last <= stage0_payload_last;
      stage0_rData_fragment_addr <= stage0_payload_fragment_addr;
      stage0_rData_fragment_id <= stage0_payload_fragment_id;
      stage0_rData_fragment_size <= stage0_payload_fragment_size;
      stage0_rData_fragment_burst <= stage0_payload_fragment_burst;
      stage0_rData_fragment_write <= stage0_payload_fragment_write;
    end
  end


endmodule

module WritebackController (
  input  wire          io_aluWrites_0_valid,
  input  wire [10:0]   io_aluWrites_0_payload_addr,
  input  wire [31:0]   io_aluWrites_0_payload_data,
  input  wire          io_valuWrites_0_valid,
  input  wire [10:0]   io_valuWrites_0_payload_addr,
  input  wire [31:0]   io_valuWrites_0_payload_data,
  input  wire          io_valuWrites_1_valid,
  input  wire [10:0]   io_valuWrites_1_payload_addr,
  input  wire [31:0]   io_valuWrites_1_payload_data,
  input  wire          io_valuWrites_2_valid,
  input  wire [10:0]   io_valuWrites_2_payload_addr,
  input  wire [31:0]   io_valuWrites_2_payload_data,
  input  wire          io_valuWrites_3_valid,
  input  wire [10:0]   io_valuWrites_3_payload_addr,
  input  wire [31:0]   io_valuWrites_3_payload_data,
  input  wire          io_valuWrites_4_valid,
  input  wire [10:0]   io_valuWrites_4_payload_addr,
  input  wire [31:0]   io_valuWrites_4_payload_data,
  input  wire          io_valuWrites_5_valid,
  input  wire [10:0]   io_valuWrites_5_payload_addr,
  input  wire [31:0]   io_valuWrites_5_payload_data,
  input  wire          io_valuWrites_6_valid,
  input  wire [10:0]   io_valuWrites_6_payload_addr,
  input  wire [31:0]   io_valuWrites_6_payload_data,
  input  wire          io_valuWrites_7_valid,
  input  wire [10:0]   io_valuWrites_7_payload_addr,
  input  wire [31:0]   io_valuWrites_7_payload_data,
  input  wire          io_loadWrites_0_valid,
  input  wire [10:0]   io_loadWrites_0_payload_addr,
  input  wire [31:0]   io_loadWrites_0_payload_data,
  input  wire          io_constWrites_0_valid,
  input  wire [10:0]   io_constWrites_0_payload_addr,
  input  wire [31:0]   io_constWrites_0_payload_data,
  input  wire          io_vloadWrites_0_valid,
  input  wire [10:0]   io_vloadWrites_0_payload_addr,
  input  wire [31:0]   io_vloadWrites_0_payload_data,
  input  wire          io_vloadWrites_1_valid,
  input  wire [10:0]   io_vloadWrites_1_payload_addr,
  input  wire [31:0]   io_vloadWrites_1_payload_data,
  input  wire          io_vloadWrites_2_valid,
  input  wire [10:0]   io_vloadWrites_2_payload_addr,
  input  wire [31:0]   io_vloadWrites_2_payload_data,
  input  wire          io_vloadWrites_3_valid,
  input  wire [10:0]   io_vloadWrites_3_payload_addr,
  input  wire [31:0]   io_vloadWrites_3_payload_data,
  input  wire          io_vloadWrites_4_valid,
  input  wire [10:0]   io_vloadWrites_4_payload_addr,
  input  wire [31:0]   io_vloadWrites_4_payload_data,
  input  wire          io_vloadWrites_5_valid,
  input  wire [10:0]   io_vloadWrites_5_payload_addr,
  input  wire [31:0]   io_vloadWrites_5_payload_data,
  input  wire          io_vloadWrites_6_valid,
  input  wire [10:0]   io_vloadWrites_6_payload_addr,
  input  wire [31:0]   io_vloadWrites_6_payload_data,
  input  wire          io_vloadWrites_7_valid,
  input  wire [10:0]   io_vloadWrites_7_payload_addr,
  input  wire [31:0]   io_vloadWrites_7_payload_data,
  input  wire          io_flowScalarWrite_valid,
  input  wire [10:0]   io_flowScalarWrite_payload_addr,
  input  wire [31:0]   io_flowScalarWrite_payload_data,
  input  wire          io_flowVectorWrites_0_valid,
  input  wire [10:0]   io_flowVectorWrites_0_payload_addr,
  input  wire [31:0]   io_flowVectorWrites_0_payload_data,
  input  wire          io_flowVectorWrites_1_valid,
  input  wire [10:0]   io_flowVectorWrites_1_payload_addr,
  input  wire [31:0]   io_flowVectorWrites_1_payload_data,
  input  wire          io_flowVectorWrites_2_valid,
  input  wire [10:0]   io_flowVectorWrites_2_payload_addr,
  input  wire [31:0]   io_flowVectorWrites_2_payload_data,
  input  wire          io_flowVectorWrites_3_valid,
  input  wire [10:0]   io_flowVectorWrites_3_payload_addr,
  input  wire [31:0]   io_flowVectorWrites_3_payload_data,
  input  wire          io_flowVectorWrites_4_valid,
  input  wire [10:0]   io_flowVectorWrites_4_payload_addr,
  input  wire [31:0]   io_flowVectorWrites_4_payload_data,
  input  wire          io_flowVectorWrites_5_valid,
  input  wire [10:0]   io_flowVectorWrites_5_payload_addr,
  input  wire [31:0]   io_flowVectorWrites_5_payload_data,
  input  wire          io_flowVectorWrites_6_valid,
  input  wire [10:0]   io_flowVectorWrites_6_payload_addr,
  input  wire [31:0]   io_flowVectorWrites_6_payload_data,
  input  wire          io_flowVectorWrites_7_valid,
  input  wire [10:0]   io_flowVectorWrites_7_payload_addr,
  input  wire [31:0]   io_flowVectorWrites_7_payload_data,
  output wire [10:0]   io_scratchWriteAddr_0,
  output wire [10:0]   io_scratchWriteAddr_1,
  output wire [10:0]   io_scratchWriteAddr_2,
  output wire [10:0]   io_scratchWriteAddr_3,
  output wire [10:0]   io_scratchWriteAddr_4,
  output wire [10:0]   io_scratchWriteAddr_5,
  output wire [10:0]   io_scratchWriteAddr_6,
  output wire [10:0]   io_scratchWriteAddr_7,
  output wire [10:0]   io_scratchWriteAddr_8,
  output wire [10:0]   io_scratchWriteAddr_9,
  output wire [10:0]   io_scratchWriteAddr_10,
  output wire [10:0]   io_scratchWriteAddr_11,
  output wire [10:0]   io_scratchWriteAddr_12,
  output wire [10:0]   io_scratchWriteAddr_13,
  output wire [10:0]   io_scratchWriteAddr_14,
  output wire [10:0]   io_scratchWriteAddr_15,
  output wire [10:0]   io_scratchWriteAddr_16,
  output wire [10:0]   io_scratchWriteAddr_17,
  output wire [10:0]   io_scratchWriteAddr_18,
  output wire [10:0]   io_scratchWriteAddr_19,
  output wire [10:0]   io_scratchWriteAddr_20,
  output wire [10:0]   io_scratchWriteAddr_21,
  output wire [10:0]   io_scratchWriteAddr_22,
  output wire [10:0]   io_scratchWriteAddr_23,
  output wire [10:0]   io_scratchWriteAddr_24,
  output wire [10:0]   io_scratchWriteAddr_25,
  output wire [10:0]   io_scratchWriteAddr_26,
  output wire [10:0]   io_scratchWriteAddr_27,
  output wire [31:0]   io_scratchWriteData_0,
  output wire [31:0]   io_scratchWriteData_1,
  output wire [31:0]   io_scratchWriteData_2,
  output wire [31:0]   io_scratchWriteData_3,
  output wire [31:0]   io_scratchWriteData_4,
  output wire [31:0]   io_scratchWriteData_5,
  output wire [31:0]   io_scratchWriteData_6,
  output wire [31:0]   io_scratchWriteData_7,
  output wire [31:0]   io_scratchWriteData_8,
  output wire [31:0]   io_scratchWriteData_9,
  output wire [31:0]   io_scratchWriteData_10,
  output wire [31:0]   io_scratchWriteData_11,
  output wire [31:0]   io_scratchWriteData_12,
  output wire [31:0]   io_scratchWriteData_13,
  output wire [31:0]   io_scratchWriteData_14,
  output wire [31:0]   io_scratchWriteData_15,
  output wire [31:0]   io_scratchWriteData_16,
  output wire [31:0]   io_scratchWriteData_17,
  output wire [31:0]   io_scratchWriteData_18,
  output wire [31:0]   io_scratchWriteData_19,
  output wire [31:0]   io_scratchWriteData_20,
  output wire [31:0]   io_scratchWriteData_21,
  output wire [31:0]   io_scratchWriteData_22,
  output wire [31:0]   io_scratchWriteData_23,
  output wire [31:0]   io_scratchWriteData_24,
  output wire [31:0]   io_scratchWriteData_25,
  output wire [31:0]   io_scratchWriteData_26,
  output wire [31:0]   io_scratchWriteData_27,
  output wire          io_scratchWriteEn_0,
  output wire          io_scratchWriteEn_1,
  output wire          io_scratchWriteEn_2,
  output wire          io_scratchWriteEn_3,
  output wire          io_scratchWriteEn_4,
  output wire          io_scratchWriteEn_5,
  output wire          io_scratchWriteEn_6,
  output wire          io_scratchWriteEn_7,
  output wire          io_scratchWriteEn_8,
  output wire          io_scratchWriteEn_9,
  output wire          io_scratchWriteEn_10,
  output wire          io_scratchWriteEn_11,
  output wire          io_scratchWriteEn_12,
  output wire          io_scratchWriteEn_13,
  output wire          io_scratchWriteEn_14,
  output wire          io_scratchWriteEn_15,
  output wire          io_scratchWriteEn_16,
  output wire          io_scratchWriteEn_17,
  output wire          io_scratchWriteEn_18,
  output wire          io_scratchWriteEn_19,
  output wire          io_scratchWriteEn_20,
  output wire          io_scratchWriteEn_21,
  output wire          io_scratchWriteEn_22,
  output wire          io_scratchWriteEn_23,
  output wire          io_scratchWriteEn_24,
  output wire          io_scratchWriteEn_25,
  output wire          io_scratchWriteEn_26,
  output wire          io_scratchWriteEn_27,
  output reg           io_wawConflict,
  input  wire          clk,
  input  wire          reset
);

  wire                when_WritebackController_l84;
  wire                when_WritebackController_l84_1;
  wire                when_WritebackController_l84_2;
  wire                when_WritebackController_l84_3;
  wire                when_WritebackController_l84_4;
  wire                when_WritebackController_l84_5;
  wire                when_WritebackController_l84_6;
  wire                when_WritebackController_l84_7;
  wire                when_WritebackController_l84_8;
  wire                when_WritebackController_l84_9;
  wire                when_WritebackController_l84_10;
  wire                when_WritebackController_l84_11;
  wire                when_WritebackController_l84_12;
  wire                when_WritebackController_l84_13;
  wire                when_WritebackController_l84_14;
  wire                when_WritebackController_l84_15;
  wire                when_WritebackController_l84_16;
  wire                when_WritebackController_l84_17;
  wire                when_WritebackController_l84_18;
  wire                when_WritebackController_l84_19;
  wire                when_WritebackController_l84_20;
  wire                when_WritebackController_l84_21;
  wire                when_WritebackController_l84_22;
  wire                when_WritebackController_l84_23;
  wire                when_WritebackController_l84_24;
  wire                when_WritebackController_l84_25;
  wire                when_WritebackController_l84_26;
  wire                when_WritebackController_l84_27;
  wire                when_WritebackController_l84_28;
  wire                when_WritebackController_l84_29;
  wire                when_WritebackController_l84_30;
  wire                when_WritebackController_l84_31;
  wire                when_WritebackController_l84_32;
  wire                when_WritebackController_l84_33;
  wire                when_WritebackController_l84_34;
  wire                when_WritebackController_l84_35;
  wire                when_WritebackController_l84_36;
  wire                when_WritebackController_l84_37;
  wire                when_WritebackController_l84_38;
  wire                when_WritebackController_l84_39;
  wire                when_WritebackController_l84_40;
  wire                when_WritebackController_l84_41;
  wire                when_WritebackController_l84_42;
  wire                when_WritebackController_l84_43;
  wire                when_WritebackController_l84_44;
  wire                when_WritebackController_l84_45;
  wire                when_WritebackController_l84_46;
  wire                when_WritebackController_l84_47;
  wire                when_WritebackController_l84_48;
  wire                when_WritebackController_l84_49;
  wire                when_WritebackController_l84_50;
  wire                when_WritebackController_l84_51;
  wire                when_WritebackController_l84_52;
  wire                when_WritebackController_l84_53;
  wire                when_WritebackController_l84_54;
  wire                when_WritebackController_l84_55;
  wire                when_WritebackController_l84_56;
  wire                when_WritebackController_l84_57;
  wire                when_WritebackController_l84_58;
  wire                when_WritebackController_l84_59;
  wire                when_WritebackController_l84_60;
  wire                when_WritebackController_l84_61;
  wire                when_WritebackController_l84_62;
  wire                when_WritebackController_l84_63;
  wire                when_WritebackController_l84_64;
  wire                when_WritebackController_l84_65;
  wire                when_WritebackController_l84_66;
  wire                when_WritebackController_l84_67;
  wire                when_WritebackController_l84_68;
  wire                when_WritebackController_l84_69;
  wire                when_WritebackController_l84_70;
  wire                when_WritebackController_l84_71;
  wire                when_WritebackController_l84_72;
  wire                when_WritebackController_l84_73;
  wire                when_WritebackController_l84_74;
  wire                when_WritebackController_l84_75;
  wire                when_WritebackController_l84_76;
  wire                when_WritebackController_l84_77;
  wire                when_WritebackController_l84_78;
  wire                when_WritebackController_l84_79;
  wire                when_WritebackController_l84_80;
  wire                when_WritebackController_l84_81;
  wire                when_WritebackController_l84_82;
  wire                when_WritebackController_l84_83;
  wire                when_WritebackController_l84_84;
  wire                when_WritebackController_l84_85;
  wire                when_WritebackController_l84_86;
  wire                when_WritebackController_l84_87;
  wire                when_WritebackController_l84_88;
  wire                when_WritebackController_l84_89;
  wire                when_WritebackController_l84_90;
  wire                when_WritebackController_l84_91;
  wire                when_WritebackController_l84_92;
  wire                when_WritebackController_l84_93;
  wire                when_WritebackController_l84_94;
  wire                when_WritebackController_l84_95;
  wire                when_WritebackController_l84_96;
  wire                when_WritebackController_l84_97;
  wire                when_WritebackController_l84_98;
  wire                when_WritebackController_l84_99;
  wire                when_WritebackController_l84_100;
  wire                when_WritebackController_l84_101;
  wire                when_WritebackController_l84_102;
  wire                when_WritebackController_l84_103;
  wire                when_WritebackController_l84_104;
  wire                when_WritebackController_l84_105;
  wire                when_WritebackController_l84_106;
  wire                when_WritebackController_l84_107;
  wire                when_WritebackController_l84_108;
  wire                when_WritebackController_l84_109;
  wire                when_WritebackController_l84_110;
  wire                when_WritebackController_l84_111;
  wire                when_WritebackController_l84_112;
  wire                when_WritebackController_l84_113;
  wire                when_WritebackController_l84_114;
  wire                when_WritebackController_l84_115;
  wire                when_WritebackController_l84_116;
  wire                when_WritebackController_l84_117;
  wire                when_WritebackController_l84_118;
  wire                when_WritebackController_l84_119;
  wire                when_WritebackController_l84_120;
  wire                when_WritebackController_l84_121;
  wire                when_WritebackController_l84_122;
  wire                when_WritebackController_l84_123;
  wire                when_WritebackController_l84_124;
  wire                when_WritebackController_l84_125;
  wire                when_WritebackController_l84_126;
  wire                when_WritebackController_l84_127;
  wire                when_WritebackController_l84_128;
  wire                when_WritebackController_l84_129;
  wire                when_WritebackController_l84_130;
  wire                when_WritebackController_l84_131;
  wire                when_WritebackController_l84_132;
  wire                when_WritebackController_l84_133;
  wire                when_WritebackController_l84_134;
  wire                when_WritebackController_l84_135;
  wire                when_WritebackController_l84_136;
  wire                when_WritebackController_l84_137;
  wire                when_WritebackController_l84_138;
  wire                when_WritebackController_l84_139;
  wire                when_WritebackController_l84_140;
  wire                when_WritebackController_l84_141;
  wire                when_WritebackController_l84_142;
  wire                when_WritebackController_l84_143;
  wire                when_WritebackController_l84_144;
  wire                when_WritebackController_l84_145;
  wire                when_WritebackController_l84_146;
  wire                when_WritebackController_l84_147;
  wire                when_WritebackController_l84_148;
  wire                when_WritebackController_l84_149;
  wire                when_WritebackController_l84_150;
  wire                when_WritebackController_l84_151;
  wire                when_WritebackController_l84_152;
  wire                when_WritebackController_l84_153;
  wire                when_WritebackController_l84_154;
  wire                when_WritebackController_l84_155;
  wire                when_WritebackController_l84_156;
  wire                when_WritebackController_l84_157;
  wire                when_WritebackController_l84_158;
  wire                when_WritebackController_l84_159;
  wire                when_WritebackController_l84_160;
  wire                when_WritebackController_l84_161;
  wire                when_WritebackController_l84_162;
  wire                when_WritebackController_l84_163;
  wire                when_WritebackController_l84_164;
  wire                when_WritebackController_l84_165;
  wire                when_WritebackController_l84_166;
  wire                when_WritebackController_l84_167;
  wire                when_WritebackController_l84_168;
  wire                when_WritebackController_l84_169;
  wire                when_WritebackController_l84_170;
  wire                when_WritebackController_l84_171;
  wire                when_WritebackController_l84_172;
  wire                when_WritebackController_l84_173;
  wire                when_WritebackController_l84_174;
  wire                when_WritebackController_l84_175;
  wire                when_WritebackController_l84_176;
  wire                when_WritebackController_l84_177;
  wire                when_WritebackController_l84_178;
  wire                when_WritebackController_l84_179;
  wire                when_WritebackController_l84_180;
  wire                when_WritebackController_l84_181;
  wire                when_WritebackController_l84_182;
  wire                when_WritebackController_l84_183;
  wire                when_WritebackController_l84_184;
  wire                when_WritebackController_l84_185;
  wire                when_WritebackController_l84_186;
  wire                when_WritebackController_l84_187;
  wire                when_WritebackController_l84_188;
  wire                when_WritebackController_l84_189;
  wire                when_WritebackController_l84_190;
  wire                when_WritebackController_l84_191;
  wire                when_WritebackController_l84_192;
  wire                when_WritebackController_l84_193;
  wire                when_WritebackController_l84_194;
  wire                when_WritebackController_l84_195;
  wire                when_WritebackController_l84_196;
  wire                when_WritebackController_l84_197;
  wire                when_WritebackController_l84_198;
  wire                when_WritebackController_l84_199;
  wire                when_WritebackController_l84_200;
  wire                when_WritebackController_l84_201;
  wire                when_WritebackController_l84_202;
  wire                when_WritebackController_l84_203;
  wire                when_WritebackController_l84_204;
  wire                when_WritebackController_l84_205;
  wire                when_WritebackController_l84_206;
  wire                when_WritebackController_l84_207;
  wire                when_WritebackController_l84_208;
  wire                when_WritebackController_l84_209;
  wire                when_WritebackController_l84_210;
  wire                when_WritebackController_l84_211;
  wire                when_WritebackController_l84_212;
  wire                when_WritebackController_l84_213;
  wire                when_WritebackController_l84_214;
  wire                when_WritebackController_l84_215;
  wire                when_WritebackController_l84_216;
  wire                when_WritebackController_l84_217;
  wire                when_WritebackController_l84_218;
  wire                when_WritebackController_l84_219;
  wire                when_WritebackController_l84_220;
  wire                when_WritebackController_l84_221;
  wire                when_WritebackController_l84_222;
  wire                when_WritebackController_l84_223;
  wire                when_WritebackController_l84_224;
  wire                when_WritebackController_l84_225;
  wire                when_WritebackController_l84_226;
  wire                when_WritebackController_l84_227;
  wire                when_WritebackController_l84_228;
  wire                when_WritebackController_l84_229;
  wire                when_WritebackController_l84_230;
  wire                when_WritebackController_l84_231;
  wire                when_WritebackController_l84_232;
  wire                when_WritebackController_l84_233;
  wire                when_WritebackController_l84_234;
  wire                when_WritebackController_l84_235;
  wire                when_WritebackController_l84_236;
  wire                when_WritebackController_l84_237;
  wire                when_WritebackController_l84_238;
  wire                when_WritebackController_l84_239;
  wire                when_WritebackController_l84_240;
  wire                when_WritebackController_l84_241;
  wire                when_WritebackController_l84_242;
  wire                when_WritebackController_l84_243;
  wire                when_WritebackController_l84_244;
  wire                when_WritebackController_l84_245;
  wire                when_WritebackController_l84_246;
  wire                when_WritebackController_l84_247;
  wire                when_WritebackController_l84_248;
  wire                when_WritebackController_l84_249;
  wire                when_WritebackController_l84_250;
  wire                when_WritebackController_l84_251;
  wire                when_WritebackController_l84_252;
  wire                when_WritebackController_l84_253;
  wire                when_WritebackController_l84_254;
  wire                when_WritebackController_l84_255;
  wire                when_WritebackController_l84_256;
  wire                when_WritebackController_l84_257;
  wire                when_WritebackController_l84_258;
  wire                when_WritebackController_l84_259;
  wire                when_WritebackController_l84_260;
  wire                when_WritebackController_l84_261;
  wire                when_WritebackController_l84_262;
  wire                when_WritebackController_l84_263;
  wire                when_WritebackController_l84_264;
  wire                when_WritebackController_l84_265;
  wire                when_WritebackController_l84_266;
  wire                when_WritebackController_l84_267;
  wire                when_WritebackController_l84_268;
  wire                when_WritebackController_l84_269;
  wire                when_WritebackController_l84_270;
  wire                when_WritebackController_l84_271;
  wire                when_WritebackController_l84_272;
  wire                when_WritebackController_l84_273;
  wire                when_WritebackController_l84_274;
  wire                when_WritebackController_l84_275;
  wire                when_WritebackController_l84_276;
  wire                when_WritebackController_l84_277;
  wire                when_WritebackController_l84_278;
  wire                when_WritebackController_l84_279;
  wire                when_WritebackController_l84_280;
  wire                when_WritebackController_l84_281;
  wire                when_WritebackController_l84_282;
  wire                when_WritebackController_l84_283;
  wire                when_WritebackController_l84_284;
  wire                when_WritebackController_l84_285;
  wire                when_WritebackController_l84_286;
  wire                when_WritebackController_l84_287;
  wire                when_WritebackController_l84_288;
  wire                when_WritebackController_l84_289;
  wire                when_WritebackController_l84_290;
  wire                when_WritebackController_l84_291;
  wire                when_WritebackController_l84_292;
  wire                when_WritebackController_l84_293;
  wire                when_WritebackController_l84_294;
  wire                when_WritebackController_l84_295;
  wire                when_WritebackController_l84_296;
  wire                when_WritebackController_l84_297;
  wire                when_WritebackController_l84_298;
  wire                when_WritebackController_l84_299;
  wire                when_WritebackController_l84_300;
  wire                when_WritebackController_l84_301;
  wire                when_WritebackController_l84_302;
  wire                when_WritebackController_l84_303;
  wire                when_WritebackController_l84_304;
  wire                when_WritebackController_l84_305;
  wire                when_WritebackController_l84_306;
  wire                when_WritebackController_l84_307;
  wire                when_WritebackController_l84_308;
  wire                when_WritebackController_l84_309;
  wire                when_WritebackController_l84_310;
  wire                when_WritebackController_l84_311;
  wire                when_WritebackController_l84_312;
  wire                when_WritebackController_l84_313;
  wire                when_WritebackController_l84_314;
  wire                when_WritebackController_l84_315;
  wire                when_WritebackController_l84_316;
  wire                when_WritebackController_l84_317;
  wire                when_WritebackController_l84_318;
  wire                when_WritebackController_l84_319;
  wire                when_WritebackController_l84_320;
  wire                when_WritebackController_l84_321;
  wire                when_WritebackController_l84_322;
  wire                when_WritebackController_l84_323;
  wire                when_WritebackController_l84_324;
  wire                when_WritebackController_l84_325;
  wire                when_WritebackController_l84_326;
  wire                when_WritebackController_l84_327;
  wire                when_WritebackController_l84_328;
  wire                when_WritebackController_l84_329;
  wire                when_WritebackController_l84_330;
  wire                when_WritebackController_l84_331;
  wire                when_WritebackController_l84_332;
  wire                when_WritebackController_l84_333;
  wire                when_WritebackController_l84_334;
  wire                when_WritebackController_l84_335;
  wire                when_WritebackController_l84_336;
  wire                when_WritebackController_l84_337;
  wire                when_WritebackController_l84_338;
  wire                when_WritebackController_l84_339;
  wire                when_WritebackController_l84_340;
  wire                when_WritebackController_l84_341;
  wire                when_WritebackController_l84_342;
  wire                when_WritebackController_l84_343;
  wire                when_WritebackController_l84_344;
  wire                when_WritebackController_l84_345;
  wire                when_WritebackController_l84_346;
  wire                when_WritebackController_l84_347;
  wire                when_WritebackController_l84_348;
  wire                when_WritebackController_l84_349;
  wire                when_WritebackController_l84_350;
  wire                when_WritebackController_l84_351;
  wire                when_WritebackController_l84_352;
  wire                when_WritebackController_l84_353;
  wire                when_WritebackController_l84_354;
  wire                when_WritebackController_l84_355;
  wire                when_WritebackController_l84_356;
  wire                when_WritebackController_l84_357;
  wire                when_WritebackController_l84_358;
  wire                when_WritebackController_l84_359;
  wire                when_WritebackController_l84_360;
  wire                when_WritebackController_l84_361;
  wire                when_WritebackController_l84_362;
  wire                when_WritebackController_l84_363;
  wire                when_WritebackController_l84_364;
  wire                when_WritebackController_l84_365;
  wire                when_WritebackController_l84_366;
  wire                when_WritebackController_l84_367;
  wire                when_WritebackController_l84_368;
  wire                when_WritebackController_l84_369;
  wire                when_WritebackController_l84_370;
  wire                when_WritebackController_l84_371;
  wire                when_WritebackController_l84_372;
  wire                when_WritebackController_l84_373;
  wire                when_WritebackController_l84_374;
  wire                when_WritebackController_l84_375;
  wire                when_WritebackController_l84_376;
  wire                when_WritebackController_l84_377;

  assign io_scratchWriteAddr_0 = io_aluWrites_0_payload_addr;
  assign io_scratchWriteData_0 = io_aluWrites_0_payload_data;
  assign io_scratchWriteEn_0 = io_aluWrites_0_valid;
  assign io_scratchWriteAddr_1 = io_valuWrites_0_payload_addr;
  assign io_scratchWriteData_1 = io_valuWrites_0_payload_data;
  assign io_scratchWriteEn_1 = io_valuWrites_0_valid;
  assign io_scratchWriteAddr_2 = io_valuWrites_1_payload_addr;
  assign io_scratchWriteData_2 = io_valuWrites_1_payload_data;
  assign io_scratchWriteEn_2 = io_valuWrites_1_valid;
  assign io_scratchWriteAddr_3 = io_valuWrites_2_payload_addr;
  assign io_scratchWriteData_3 = io_valuWrites_2_payload_data;
  assign io_scratchWriteEn_3 = io_valuWrites_2_valid;
  assign io_scratchWriteAddr_4 = io_valuWrites_3_payload_addr;
  assign io_scratchWriteData_4 = io_valuWrites_3_payload_data;
  assign io_scratchWriteEn_4 = io_valuWrites_3_valid;
  assign io_scratchWriteAddr_5 = io_valuWrites_4_payload_addr;
  assign io_scratchWriteData_5 = io_valuWrites_4_payload_data;
  assign io_scratchWriteEn_5 = io_valuWrites_4_valid;
  assign io_scratchWriteAddr_6 = io_valuWrites_5_payload_addr;
  assign io_scratchWriteData_6 = io_valuWrites_5_payload_data;
  assign io_scratchWriteEn_6 = io_valuWrites_5_valid;
  assign io_scratchWriteAddr_7 = io_valuWrites_6_payload_addr;
  assign io_scratchWriteData_7 = io_valuWrites_6_payload_data;
  assign io_scratchWriteEn_7 = io_valuWrites_6_valid;
  assign io_scratchWriteAddr_8 = io_valuWrites_7_payload_addr;
  assign io_scratchWriteData_8 = io_valuWrites_7_payload_data;
  assign io_scratchWriteEn_8 = io_valuWrites_7_valid;
  assign io_scratchWriteAddr_9 = io_loadWrites_0_payload_addr;
  assign io_scratchWriteData_9 = io_loadWrites_0_payload_data;
  assign io_scratchWriteEn_9 = io_loadWrites_0_valid;
  assign io_scratchWriteAddr_10 = io_constWrites_0_payload_addr;
  assign io_scratchWriteData_10 = io_constWrites_0_payload_data;
  assign io_scratchWriteEn_10 = io_constWrites_0_valid;
  assign io_scratchWriteAddr_11 = io_vloadWrites_0_payload_addr;
  assign io_scratchWriteData_11 = io_vloadWrites_0_payload_data;
  assign io_scratchWriteEn_11 = io_vloadWrites_0_valid;
  assign io_scratchWriteAddr_12 = io_vloadWrites_1_payload_addr;
  assign io_scratchWriteData_12 = io_vloadWrites_1_payload_data;
  assign io_scratchWriteEn_12 = io_vloadWrites_1_valid;
  assign io_scratchWriteAddr_13 = io_vloadWrites_2_payload_addr;
  assign io_scratchWriteData_13 = io_vloadWrites_2_payload_data;
  assign io_scratchWriteEn_13 = io_vloadWrites_2_valid;
  assign io_scratchWriteAddr_14 = io_vloadWrites_3_payload_addr;
  assign io_scratchWriteData_14 = io_vloadWrites_3_payload_data;
  assign io_scratchWriteEn_14 = io_vloadWrites_3_valid;
  assign io_scratchWriteAddr_15 = io_vloadWrites_4_payload_addr;
  assign io_scratchWriteData_15 = io_vloadWrites_4_payload_data;
  assign io_scratchWriteEn_15 = io_vloadWrites_4_valid;
  assign io_scratchWriteAddr_16 = io_vloadWrites_5_payload_addr;
  assign io_scratchWriteData_16 = io_vloadWrites_5_payload_data;
  assign io_scratchWriteEn_16 = io_vloadWrites_5_valid;
  assign io_scratchWriteAddr_17 = io_vloadWrites_6_payload_addr;
  assign io_scratchWriteData_17 = io_vloadWrites_6_payload_data;
  assign io_scratchWriteEn_17 = io_vloadWrites_6_valid;
  assign io_scratchWriteAddr_18 = io_vloadWrites_7_payload_addr;
  assign io_scratchWriteData_18 = io_vloadWrites_7_payload_data;
  assign io_scratchWriteEn_18 = io_vloadWrites_7_valid;
  assign io_scratchWriteAddr_19 = io_flowScalarWrite_payload_addr;
  assign io_scratchWriteData_19 = io_flowScalarWrite_payload_data;
  assign io_scratchWriteEn_19 = io_flowScalarWrite_valid;
  assign io_scratchWriteAddr_20 = io_flowVectorWrites_0_payload_addr;
  assign io_scratchWriteData_20 = io_flowVectorWrites_0_payload_data;
  assign io_scratchWriteEn_20 = io_flowVectorWrites_0_valid;
  assign io_scratchWriteAddr_21 = io_flowVectorWrites_1_payload_addr;
  assign io_scratchWriteData_21 = io_flowVectorWrites_1_payload_data;
  assign io_scratchWriteEn_21 = io_flowVectorWrites_1_valid;
  assign io_scratchWriteAddr_22 = io_flowVectorWrites_2_payload_addr;
  assign io_scratchWriteData_22 = io_flowVectorWrites_2_payload_data;
  assign io_scratchWriteEn_22 = io_flowVectorWrites_2_valid;
  assign io_scratchWriteAddr_23 = io_flowVectorWrites_3_payload_addr;
  assign io_scratchWriteData_23 = io_flowVectorWrites_3_payload_data;
  assign io_scratchWriteEn_23 = io_flowVectorWrites_3_valid;
  assign io_scratchWriteAddr_24 = io_flowVectorWrites_4_payload_addr;
  assign io_scratchWriteData_24 = io_flowVectorWrites_4_payload_data;
  assign io_scratchWriteEn_24 = io_flowVectorWrites_4_valid;
  assign io_scratchWriteAddr_25 = io_flowVectorWrites_5_payload_addr;
  assign io_scratchWriteData_25 = io_flowVectorWrites_5_payload_data;
  assign io_scratchWriteEn_25 = io_flowVectorWrites_5_valid;
  assign io_scratchWriteAddr_26 = io_flowVectorWrites_6_payload_addr;
  assign io_scratchWriteData_26 = io_flowVectorWrites_6_payload_data;
  assign io_scratchWriteEn_26 = io_flowVectorWrites_6_valid;
  assign io_scratchWriteAddr_27 = io_flowVectorWrites_7_payload_addr;
  assign io_scratchWriteData_27 = io_flowVectorWrites_7_payload_data;
  assign io_scratchWriteEn_27 = io_flowVectorWrites_7_valid;
  always @(*) begin
    io_wawConflict = 1'b0;
    if(when_WritebackController_l84) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_1) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_2) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_3) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_4) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_5) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_6) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_7) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_8) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_9) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_10) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_11) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_12) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_13) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_14) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_15) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_16) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_17) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_18) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_19) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_20) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_21) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_22) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_23) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_24) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_25) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_26) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_27) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_28) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_29) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_30) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_31) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_32) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_33) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_34) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_35) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_36) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_37) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_38) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_39) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_40) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_41) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_42) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_43) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_44) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_45) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_46) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_47) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_48) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_49) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_50) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_51) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_52) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_53) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_54) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_55) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_56) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_57) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_58) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_59) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_60) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_61) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_62) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_63) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_64) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_65) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_66) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_67) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_68) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_69) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_70) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_71) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_72) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_73) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_74) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_75) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_76) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_77) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_78) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_79) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_80) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_81) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_82) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_83) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_84) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_85) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_86) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_87) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_88) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_89) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_90) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_91) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_92) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_93) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_94) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_95) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_96) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_97) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_98) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_99) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_100) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_101) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_102) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_103) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_104) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_105) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_106) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_107) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_108) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_109) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_110) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_111) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_112) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_113) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_114) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_115) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_116) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_117) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_118) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_119) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_120) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_121) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_122) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_123) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_124) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_125) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_126) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_127) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_128) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_129) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_130) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_131) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_132) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_133) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_134) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_135) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_136) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_137) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_138) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_139) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_140) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_141) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_142) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_143) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_144) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_145) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_146) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_147) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_148) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_149) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_150) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_151) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_152) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_153) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_154) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_155) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_156) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_157) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_158) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_159) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_160) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_161) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_162) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_163) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_164) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_165) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_166) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_167) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_168) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_169) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_170) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_171) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_172) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_173) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_174) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_175) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_176) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_177) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_178) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_179) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_180) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_181) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_182) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_183) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_184) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_185) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_186) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_187) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_188) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_189) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_190) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_191) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_192) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_193) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_194) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_195) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_196) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_197) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_198) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_199) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_200) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_201) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_202) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_203) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_204) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_205) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_206) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_207) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_208) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_209) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_210) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_211) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_212) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_213) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_214) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_215) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_216) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_217) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_218) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_219) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_220) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_221) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_222) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_223) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_224) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_225) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_226) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_227) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_228) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_229) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_230) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_231) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_232) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_233) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_234) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_235) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_236) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_237) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_238) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_239) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_240) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_241) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_242) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_243) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_244) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_245) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_246) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_247) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_248) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_249) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_250) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_251) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_252) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_253) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_254) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_255) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_256) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_257) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_258) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_259) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_260) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_261) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_262) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_263) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_264) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_265) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_266) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_267) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_268) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_269) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_270) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_271) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_272) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_273) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_274) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_275) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_276) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_277) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_278) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_279) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_280) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_281) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_282) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_283) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_284) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_285) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_286) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_287) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_288) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_289) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_290) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_291) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_292) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_293) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_294) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_295) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_296) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_297) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_298) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_299) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_300) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_301) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_302) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_303) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_304) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_305) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_306) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_307) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_308) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_309) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_310) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_311) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_312) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_313) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_314) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_315) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_316) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_317) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_318) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_319) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_320) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_321) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_322) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_323) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_324) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_325) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_326) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_327) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_328) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_329) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_330) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_331) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_332) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_333) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_334) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_335) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_336) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_337) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_338) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_339) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_340) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_341) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_342) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_343) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_344) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_345) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_346) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_347) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_348) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_349) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_350) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_351) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_352) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_353) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_354) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_355) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_356) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_357) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_358) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_359) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_360) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_361) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_362) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_363) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_364) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_365) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_366) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_367) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_368) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_369) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_370) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_371) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_372) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_373) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_374) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_375) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_376) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l84_377) begin
      io_wawConflict = 1'b1;
    end
  end

  assign when_WritebackController_l84 = ((io_aluWrites_0_valid && io_valuWrites_0_valid) && (io_aluWrites_0_payload_addr == io_valuWrites_0_payload_addr));
  assign when_WritebackController_l84_1 = ((io_aluWrites_0_valid && io_valuWrites_1_valid) && (io_aluWrites_0_payload_addr == io_valuWrites_1_payload_addr));
  assign when_WritebackController_l84_2 = ((io_aluWrites_0_valid && io_valuWrites_2_valid) && (io_aluWrites_0_payload_addr == io_valuWrites_2_payload_addr));
  assign when_WritebackController_l84_3 = ((io_aluWrites_0_valid && io_valuWrites_3_valid) && (io_aluWrites_0_payload_addr == io_valuWrites_3_payload_addr));
  assign when_WritebackController_l84_4 = ((io_aluWrites_0_valid && io_valuWrites_4_valid) && (io_aluWrites_0_payload_addr == io_valuWrites_4_payload_addr));
  assign when_WritebackController_l84_5 = ((io_aluWrites_0_valid && io_valuWrites_5_valid) && (io_aluWrites_0_payload_addr == io_valuWrites_5_payload_addr));
  assign when_WritebackController_l84_6 = ((io_aluWrites_0_valid && io_valuWrites_6_valid) && (io_aluWrites_0_payload_addr == io_valuWrites_6_payload_addr));
  assign when_WritebackController_l84_7 = ((io_aluWrites_0_valid && io_valuWrites_7_valid) && (io_aluWrites_0_payload_addr == io_valuWrites_7_payload_addr));
  assign when_WritebackController_l84_8 = ((io_aluWrites_0_valid && io_loadWrites_0_valid) && (io_aluWrites_0_payload_addr == io_loadWrites_0_payload_addr));
  assign when_WritebackController_l84_9 = ((io_aluWrites_0_valid && io_constWrites_0_valid) && (io_aluWrites_0_payload_addr == io_constWrites_0_payload_addr));
  assign when_WritebackController_l84_10 = ((io_aluWrites_0_valid && io_vloadWrites_0_valid) && (io_aluWrites_0_payload_addr == io_vloadWrites_0_payload_addr));
  assign when_WritebackController_l84_11 = ((io_aluWrites_0_valid && io_vloadWrites_1_valid) && (io_aluWrites_0_payload_addr == io_vloadWrites_1_payload_addr));
  assign when_WritebackController_l84_12 = ((io_aluWrites_0_valid && io_vloadWrites_2_valid) && (io_aluWrites_0_payload_addr == io_vloadWrites_2_payload_addr));
  assign when_WritebackController_l84_13 = ((io_aluWrites_0_valid && io_vloadWrites_3_valid) && (io_aluWrites_0_payload_addr == io_vloadWrites_3_payload_addr));
  assign when_WritebackController_l84_14 = ((io_aluWrites_0_valid && io_vloadWrites_4_valid) && (io_aluWrites_0_payload_addr == io_vloadWrites_4_payload_addr));
  assign when_WritebackController_l84_15 = ((io_aluWrites_0_valid && io_vloadWrites_5_valid) && (io_aluWrites_0_payload_addr == io_vloadWrites_5_payload_addr));
  assign when_WritebackController_l84_16 = ((io_aluWrites_0_valid && io_vloadWrites_6_valid) && (io_aluWrites_0_payload_addr == io_vloadWrites_6_payload_addr));
  assign when_WritebackController_l84_17 = ((io_aluWrites_0_valid && io_vloadWrites_7_valid) && (io_aluWrites_0_payload_addr == io_vloadWrites_7_payload_addr));
  assign when_WritebackController_l84_18 = ((io_aluWrites_0_valid && io_flowScalarWrite_valid) && (io_aluWrites_0_payload_addr == io_flowScalarWrite_payload_addr));
  assign when_WritebackController_l84_19 = ((io_aluWrites_0_valid && io_flowVectorWrites_0_valid) && (io_aluWrites_0_payload_addr == io_flowVectorWrites_0_payload_addr));
  assign when_WritebackController_l84_20 = ((io_aluWrites_0_valid && io_flowVectorWrites_1_valid) && (io_aluWrites_0_payload_addr == io_flowVectorWrites_1_payload_addr));
  assign when_WritebackController_l84_21 = ((io_aluWrites_0_valid && io_flowVectorWrites_2_valid) && (io_aluWrites_0_payload_addr == io_flowVectorWrites_2_payload_addr));
  assign when_WritebackController_l84_22 = ((io_aluWrites_0_valid && io_flowVectorWrites_3_valid) && (io_aluWrites_0_payload_addr == io_flowVectorWrites_3_payload_addr));
  assign when_WritebackController_l84_23 = ((io_aluWrites_0_valid && io_flowVectorWrites_4_valid) && (io_aluWrites_0_payload_addr == io_flowVectorWrites_4_payload_addr));
  assign when_WritebackController_l84_24 = ((io_aluWrites_0_valid && io_flowVectorWrites_5_valid) && (io_aluWrites_0_payload_addr == io_flowVectorWrites_5_payload_addr));
  assign when_WritebackController_l84_25 = ((io_aluWrites_0_valid && io_flowVectorWrites_6_valid) && (io_aluWrites_0_payload_addr == io_flowVectorWrites_6_payload_addr));
  assign when_WritebackController_l84_26 = ((io_aluWrites_0_valid && io_flowVectorWrites_7_valid) && (io_aluWrites_0_payload_addr == io_flowVectorWrites_7_payload_addr));
  assign when_WritebackController_l84_27 = ((io_valuWrites_0_valid && io_valuWrites_1_valid) && (io_valuWrites_0_payload_addr == io_valuWrites_1_payload_addr));
  assign when_WritebackController_l84_28 = ((io_valuWrites_0_valid && io_valuWrites_2_valid) && (io_valuWrites_0_payload_addr == io_valuWrites_2_payload_addr));
  assign when_WritebackController_l84_29 = ((io_valuWrites_0_valid && io_valuWrites_3_valid) && (io_valuWrites_0_payload_addr == io_valuWrites_3_payload_addr));
  assign when_WritebackController_l84_30 = ((io_valuWrites_0_valid && io_valuWrites_4_valid) && (io_valuWrites_0_payload_addr == io_valuWrites_4_payload_addr));
  assign when_WritebackController_l84_31 = ((io_valuWrites_0_valid && io_valuWrites_5_valid) && (io_valuWrites_0_payload_addr == io_valuWrites_5_payload_addr));
  assign when_WritebackController_l84_32 = ((io_valuWrites_0_valid && io_valuWrites_6_valid) && (io_valuWrites_0_payload_addr == io_valuWrites_6_payload_addr));
  assign when_WritebackController_l84_33 = ((io_valuWrites_0_valid && io_valuWrites_7_valid) && (io_valuWrites_0_payload_addr == io_valuWrites_7_payload_addr));
  assign when_WritebackController_l84_34 = ((io_valuWrites_0_valid && io_loadWrites_0_valid) && (io_valuWrites_0_payload_addr == io_loadWrites_0_payload_addr));
  assign when_WritebackController_l84_35 = ((io_valuWrites_0_valid && io_constWrites_0_valid) && (io_valuWrites_0_payload_addr == io_constWrites_0_payload_addr));
  assign when_WritebackController_l84_36 = ((io_valuWrites_0_valid && io_vloadWrites_0_valid) && (io_valuWrites_0_payload_addr == io_vloadWrites_0_payload_addr));
  assign when_WritebackController_l84_37 = ((io_valuWrites_0_valid && io_vloadWrites_1_valid) && (io_valuWrites_0_payload_addr == io_vloadWrites_1_payload_addr));
  assign when_WritebackController_l84_38 = ((io_valuWrites_0_valid && io_vloadWrites_2_valid) && (io_valuWrites_0_payload_addr == io_vloadWrites_2_payload_addr));
  assign when_WritebackController_l84_39 = ((io_valuWrites_0_valid && io_vloadWrites_3_valid) && (io_valuWrites_0_payload_addr == io_vloadWrites_3_payload_addr));
  assign when_WritebackController_l84_40 = ((io_valuWrites_0_valid && io_vloadWrites_4_valid) && (io_valuWrites_0_payload_addr == io_vloadWrites_4_payload_addr));
  assign when_WritebackController_l84_41 = ((io_valuWrites_0_valid && io_vloadWrites_5_valid) && (io_valuWrites_0_payload_addr == io_vloadWrites_5_payload_addr));
  assign when_WritebackController_l84_42 = ((io_valuWrites_0_valid && io_vloadWrites_6_valid) && (io_valuWrites_0_payload_addr == io_vloadWrites_6_payload_addr));
  assign when_WritebackController_l84_43 = ((io_valuWrites_0_valid && io_vloadWrites_7_valid) && (io_valuWrites_0_payload_addr == io_vloadWrites_7_payload_addr));
  assign when_WritebackController_l84_44 = ((io_valuWrites_0_valid && io_flowScalarWrite_valid) && (io_valuWrites_0_payload_addr == io_flowScalarWrite_payload_addr));
  assign when_WritebackController_l84_45 = ((io_valuWrites_0_valid && io_flowVectorWrites_0_valid) && (io_valuWrites_0_payload_addr == io_flowVectorWrites_0_payload_addr));
  assign when_WritebackController_l84_46 = ((io_valuWrites_0_valid && io_flowVectorWrites_1_valid) && (io_valuWrites_0_payload_addr == io_flowVectorWrites_1_payload_addr));
  assign when_WritebackController_l84_47 = ((io_valuWrites_0_valid && io_flowVectorWrites_2_valid) && (io_valuWrites_0_payload_addr == io_flowVectorWrites_2_payload_addr));
  assign when_WritebackController_l84_48 = ((io_valuWrites_0_valid && io_flowVectorWrites_3_valid) && (io_valuWrites_0_payload_addr == io_flowVectorWrites_3_payload_addr));
  assign when_WritebackController_l84_49 = ((io_valuWrites_0_valid && io_flowVectorWrites_4_valid) && (io_valuWrites_0_payload_addr == io_flowVectorWrites_4_payload_addr));
  assign when_WritebackController_l84_50 = ((io_valuWrites_0_valid && io_flowVectorWrites_5_valid) && (io_valuWrites_0_payload_addr == io_flowVectorWrites_5_payload_addr));
  assign when_WritebackController_l84_51 = ((io_valuWrites_0_valid && io_flowVectorWrites_6_valid) && (io_valuWrites_0_payload_addr == io_flowVectorWrites_6_payload_addr));
  assign when_WritebackController_l84_52 = ((io_valuWrites_0_valid && io_flowVectorWrites_7_valid) && (io_valuWrites_0_payload_addr == io_flowVectorWrites_7_payload_addr));
  assign when_WritebackController_l84_53 = ((io_valuWrites_1_valid && io_valuWrites_2_valid) && (io_valuWrites_1_payload_addr == io_valuWrites_2_payload_addr));
  assign when_WritebackController_l84_54 = ((io_valuWrites_1_valid && io_valuWrites_3_valid) && (io_valuWrites_1_payload_addr == io_valuWrites_3_payload_addr));
  assign when_WritebackController_l84_55 = ((io_valuWrites_1_valid && io_valuWrites_4_valid) && (io_valuWrites_1_payload_addr == io_valuWrites_4_payload_addr));
  assign when_WritebackController_l84_56 = ((io_valuWrites_1_valid && io_valuWrites_5_valid) && (io_valuWrites_1_payload_addr == io_valuWrites_5_payload_addr));
  assign when_WritebackController_l84_57 = ((io_valuWrites_1_valid && io_valuWrites_6_valid) && (io_valuWrites_1_payload_addr == io_valuWrites_6_payload_addr));
  assign when_WritebackController_l84_58 = ((io_valuWrites_1_valid && io_valuWrites_7_valid) && (io_valuWrites_1_payload_addr == io_valuWrites_7_payload_addr));
  assign when_WritebackController_l84_59 = ((io_valuWrites_1_valid && io_loadWrites_0_valid) && (io_valuWrites_1_payload_addr == io_loadWrites_0_payload_addr));
  assign when_WritebackController_l84_60 = ((io_valuWrites_1_valid && io_constWrites_0_valid) && (io_valuWrites_1_payload_addr == io_constWrites_0_payload_addr));
  assign when_WritebackController_l84_61 = ((io_valuWrites_1_valid && io_vloadWrites_0_valid) && (io_valuWrites_1_payload_addr == io_vloadWrites_0_payload_addr));
  assign when_WritebackController_l84_62 = ((io_valuWrites_1_valid && io_vloadWrites_1_valid) && (io_valuWrites_1_payload_addr == io_vloadWrites_1_payload_addr));
  assign when_WritebackController_l84_63 = ((io_valuWrites_1_valid && io_vloadWrites_2_valid) && (io_valuWrites_1_payload_addr == io_vloadWrites_2_payload_addr));
  assign when_WritebackController_l84_64 = ((io_valuWrites_1_valid && io_vloadWrites_3_valid) && (io_valuWrites_1_payload_addr == io_vloadWrites_3_payload_addr));
  assign when_WritebackController_l84_65 = ((io_valuWrites_1_valid && io_vloadWrites_4_valid) && (io_valuWrites_1_payload_addr == io_vloadWrites_4_payload_addr));
  assign when_WritebackController_l84_66 = ((io_valuWrites_1_valid && io_vloadWrites_5_valid) && (io_valuWrites_1_payload_addr == io_vloadWrites_5_payload_addr));
  assign when_WritebackController_l84_67 = ((io_valuWrites_1_valid && io_vloadWrites_6_valid) && (io_valuWrites_1_payload_addr == io_vloadWrites_6_payload_addr));
  assign when_WritebackController_l84_68 = ((io_valuWrites_1_valid && io_vloadWrites_7_valid) && (io_valuWrites_1_payload_addr == io_vloadWrites_7_payload_addr));
  assign when_WritebackController_l84_69 = ((io_valuWrites_1_valid && io_flowScalarWrite_valid) && (io_valuWrites_1_payload_addr == io_flowScalarWrite_payload_addr));
  assign when_WritebackController_l84_70 = ((io_valuWrites_1_valid && io_flowVectorWrites_0_valid) && (io_valuWrites_1_payload_addr == io_flowVectorWrites_0_payload_addr));
  assign when_WritebackController_l84_71 = ((io_valuWrites_1_valid && io_flowVectorWrites_1_valid) && (io_valuWrites_1_payload_addr == io_flowVectorWrites_1_payload_addr));
  assign when_WritebackController_l84_72 = ((io_valuWrites_1_valid && io_flowVectorWrites_2_valid) && (io_valuWrites_1_payload_addr == io_flowVectorWrites_2_payload_addr));
  assign when_WritebackController_l84_73 = ((io_valuWrites_1_valid && io_flowVectorWrites_3_valid) && (io_valuWrites_1_payload_addr == io_flowVectorWrites_3_payload_addr));
  assign when_WritebackController_l84_74 = ((io_valuWrites_1_valid && io_flowVectorWrites_4_valid) && (io_valuWrites_1_payload_addr == io_flowVectorWrites_4_payload_addr));
  assign when_WritebackController_l84_75 = ((io_valuWrites_1_valid && io_flowVectorWrites_5_valid) && (io_valuWrites_1_payload_addr == io_flowVectorWrites_5_payload_addr));
  assign when_WritebackController_l84_76 = ((io_valuWrites_1_valid && io_flowVectorWrites_6_valid) && (io_valuWrites_1_payload_addr == io_flowVectorWrites_6_payload_addr));
  assign when_WritebackController_l84_77 = ((io_valuWrites_1_valid && io_flowVectorWrites_7_valid) && (io_valuWrites_1_payload_addr == io_flowVectorWrites_7_payload_addr));
  assign when_WritebackController_l84_78 = ((io_valuWrites_2_valid && io_valuWrites_3_valid) && (io_valuWrites_2_payload_addr == io_valuWrites_3_payload_addr));
  assign when_WritebackController_l84_79 = ((io_valuWrites_2_valid && io_valuWrites_4_valid) && (io_valuWrites_2_payload_addr == io_valuWrites_4_payload_addr));
  assign when_WritebackController_l84_80 = ((io_valuWrites_2_valid && io_valuWrites_5_valid) && (io_valuWrites_2_payload_addr == io_valuWrites_5_payload_addr));
  assign when_WritebackController_l84_81 = ((io_valuWrites_2_valid && io_valuWrites_6_valid) && (io_valuWrites_2_payload_addr == io_valuWrites_6_payload_addr));
  assign when_WritebackController_l84_82 = ((io_valuWrites_2_valid && io_valuWrites_7_valid) && (io_valuWrites_2_payload_addr == io_valuWrites_7_payload_addr));
  assign when_WritebackController_l84_83 = ((io_valuWrites_2_valid && io_loadWrites_0_valid) && (io_valuWrites_2_payload_addr == io_loadWrites_0_payload_addr));
  assign when_WritebackController_l84_84 = ((io_valuWrites_2_valid && io_constWrites_0_valid) && (io_valuWrites_2_payload_addr == io_constWrites_0_payload_addr));
  assign when_WritebackController_l84_85 = ((io_valuWrites_2_valid && io_vloadWrites_0_valid) && (io_valuWrites_2_payload_addr == io_vloadWrites_0_payload_addr));
  assign when_WritebackController_l84_86 = ((io_valuWrites_2_valid && io_vloadWrites_1_valid) && (io_valuWrites_2_payload_addr == io_vloadWrites_1_payload_addr));
  assign when_WritebackController_l84_87 = ((io_valuWrites_2_valid && io_vloadWrites_2_valid) && (io_valuWrites_2_payload_addr == io_vloadWrites_2_payload_addr));
  assign when_WritebackController_l84_88 = ((io_valuWrites_2_valid && io_vloadWrites_3_valid) && (io_valuWrites_2_payload_addr == io_vloadWrites_3_payload_addr));
  assign when_WritebackController_l84_89 = ((io_valuWrites_2_valid && io_vloadWrites_4_valid) && (io_valuWrites_2_payload_addr == io_vloadWrites_4_payload_addr));
  assign when_WritebackController_l84_90 = ((io_valuWrites_2_valid && io_vloadWrites_5_valid) && (io_valuWrites_2_payload_addr == io_vloadWrites_5_payload_addr));
  assign when_WritebackController_l84_91 = ((io_valuWrites_2_valid && io_vloadWrites_6_valid) && (io_valuWrites_2_payload_addr == io_vloadWrites_6_payload_addr));
  assign when_WritebackController_l84_92 = ((io_valuWrites_2_valid && io_vloadWrites_7_valid) && (io_valuWrites_2_payload_addr == io_vloadWrites_7_payload_addr));
  assign when_WritebackController_l84_93 = ((io_valuWrites_2_valid && io_flowScalarWrite_valid) && (io_valuWrites_2_payload_addr == io_flowScalarWrite_payload_addr));
  assign when_WritebackController_l84_94 = ((io_valuWrites_2_valid && io_flowVectorWrites_0_valid) && (io_valuWrites_2_payload_addr == io_flowVectorWrites_0_payload_addr));
  assign when_WritebackController_l84_95 = ((io_valuWrites_2_valid && io_flowVectorWrites_1_valid) && (io_valuWrites_2_payload_addr == io_flowVectorWrites_1_payload_addr));
  assign when_WritebackController_l84_96 = ((io_valuWrites_2_valid && io_flowVectorWrites_2_valid) && (io_valuWrites_2_payload_addr == io_flowVectorWrites_2_payload_addr));
  assign when_WritebackController_l84_97 = ((io_valuWrites_2_valid && io_flowVectorWrites_3_valid) && (io_valuWrites_2_payload_addr == io_flowVectorWrites_3_payload_addr));
  assign when_WritebackController_l84_98 = ((io_valuWrites_2_valid && io_flowVectorWrites_4_valid) && (io_valuWrites_2_payload_addr == io_flowVectorWrites_4_payload_addr));
  assign when_WritebackController_l84_99 = ((io_valuWrites_2_valid && io_flowVectorWrites_5_valid) && (io_valuWrites_2_payload_addr == io_flowVectorWrites_5_payload_addr));
  assign when_WritebackController_l84_100 = ((io_valuWrites_2_valid && io_flowVectorWrites_6_valid) && (io_valuWrites_2_payload_addr == io_flowVectorWrites_6_payload_addr));
  assign when_WritebackController_l84_101 = ((io_valuWrites_2_valid && io_flowVectorWrites_7_valid) && (io_valuWrites_2_payload_addr == io_flowVectorWrites_7_payload_addr));
  assign when_WritebackController_l84_102 = ((io_valuWrites_3_valid && io_valuWrites_4_valid) && (io_valuWrites_3_payload_addr == io_valuWrites_4_payload_addr));
  assign when_WritebackController_l84_103 = ((io_valuWrites_3_valid && io_valuWrites_5_valid) && (io_valuWrites_3_payload_addr == io_valuWrites_5_payload_addr));
  assign when_WritebackController_l84_104 = ((io_valuWrites_3_valid && io_valuWrites_6_valid) && (io_valuWrites_3_payload_addr == io_valuWrites_6_payload_addr));
  assign when_WritebackController_l84_105 = ((io_valuWrites_3_valid && io_valuWrites_7_valid) && (io_valuWrites_3_payload_addr == io_valuWrites_7_payload_addr));
  assign when_WritebackController_l84_106 = ((io_valuWrites_3_valid && io_loadWrites_0_valid) && (io_valuWrites_3_payload_addr == io_loadWrites_0_payload_addr));
  assign when_WritebackController_l84_107 = ((io_valuWrites_3_valid && io_constWrites_0_valid) && (io_valuWrites_3_payload_addr == io_constWrites_0_payload_addr));
  assign when_WritebackController_l84_108 = ((io_valuWrites_3_valid && io_vloadWrites_0_valid) && (io_valuWrites_3_payload_addr == io_vloadWrites_0_payload_addr));
  assign when_WritebackController_l84_109 = ((io_valuWrites_3_valid && io_vloadWrites_1_valid) && (io_valuWrites_3_payload_addr == io_vloadWrites_1_payload_addr));
  assign when_WritebackController_l84_110 = ((io_valuWrites_3_valid && io_vloadWrites_2_valid) && (io_valuWrites_3_payload_addr == io_vloadWrites_2_payload_addr));
  assign when_WritebackController_l84_111 = ((io_valuWrites_3_valid && io_vloadWrites_3_valid) && (io_valuWrites_3_payload_addr == io_vloadWrites_3_payload_addr));
  assign when_WritebackController_l84_112 = ((io_valuWrites_3_valid && io_vloadWrites_4_valid) && (io_valuWrites_3_payload_addr == io_vloadWrites_4_payload_addr));
  assign when_WritebackController_l84_113 = ((io_valuWrites_3_valid && io_vloadWrites_5_valid) && (io_valuWrites_3_payload_addr == io_vloadWrites_5_payload_addr));
  assign when_WritebackController_l84_114 = ((io_valuWrites_3_valid && io_vloadWrites_6_valid) && (io_valuWrites_3_payload_addr == io_vloadWrites_6_payload_addr));
  assign when_WritebackController_l84_115 = ((io_valuWrites_3_valid && io_vloadWrites_7_valid) && (io_valuWrites_3_payload_addr == io_vloadWrites_7_payload_addr));
  assign when_WritebackController_l84_116 = ((io_valuWrites_3_valid && io_flowScalarWrite_valid) && (io_valuWrites_3_payload_addr == io_flowScalarWrite_payload_addr));
  assign when_WritebackController_l84_117 = ((io_valuWrites_3_valid && io_flowVectorWrites_0_valid) && (io_valuWrites_3_payload_addr == io_flowVectorWrites_0_payload_addr));
  assign when_WritebackController_l84_118 = ((io_valuWrites_3_valid && io_flowVectorWrites_1_valid) && (io_valuWrites_3_payload_addr == io_flowVectorWrites_1_payload_addr));
  assign when_WritebackController_l84_119 = ((io_valuWrites_3_valid && io_flowVectorWrites_2_valid) && (io_valuWrites_3_payload_addr == io_flowVectorWrites_2_payload_addr));
  assign when_WritebackController_l84_120 = ((io_valuWrites_3_valid && io_flowVectorWrites_3_valid) && (io_valuWrites_3_payload_addr == io_flowVectorWrites_3_payload_addr));
  assign when_WritebackController_l84_121 = ((io_valuWrites_3_valid && io_flowVectorWrites_4_valid) && (io_valuWrites_3_payload_addr == io_flowVectorWrites_4_payload_addr));
  assign when_WritebackController_l84_122 = ((io_valuWrites_3_valid && io_flowVectorWrites_5_valid) && (io_valuWrites_3_payload_addr == io_flowVectorWrites_5_payload_addr));
  assign when_WritebackController_l84_123 = ((io_valuWrites_3_valid && io_flowVectorWrites_6_valid) && (io_valuWrites_3_payload_addr == io_flowVectorWrites_6_payload_addr));
  assign when_WritebackController_l84_124 = ((io_valuWrites_3_valid && io_flowVectorWrites_7_valid) && (io_valuWrites_3_payload_addr == io_flowVectorWrites_7_payload_addr));
  assign when_WritebackController_l84_125 = ((io_valuWrites_4_valid && io_valuWrites_5_valid) && (io_valuWrites_4_payload_addr == io_valuWrites_5_payload_addr));
  assign when_WritebackController_l84_126 = ((io_valuWrites_4_valid && io_valuWrites_6_valid) && (io_valuWrites_4_payload_addr == io_valuWrites_6_payload_addr));
  assign when_WritebackController_l84_127 = ((io_valuWrites_4_valid && io_valuWrites_7_valid) && (io_valuWrites_4_payload_addr == io_valuWrites_7_payload_addr));
  assign when_WritebackController_l84_128 = ((io_valuWrites_4_valid && io_loadWrites_0_valid) && (io_valuWrites_4_payload_addr == io_loadWrites_0_payload_addr));
  assign when_WritebackController_l84_129 = ((io_valuWrites_4_valid && io_constWrites_0_valid) && (io_valuWrites_4_payload_addr == io_constWrites_0_payload_addr));
  assign when_WritebackController_l84_130 = ((io_valuWrites_4_valid && io_vloadWrites_0_valid) && (io_valuWrites_4_payload_addr == io_vloadWrites_0_payload_addr));
  assign when_WritebackController_l84_131 = ((io_valuWrites_4_valid && io_vloadWrites_1_valid) && (io_valuWrites_4_payload_addr == io_vloadWrites_1_payload_addr));
  assign when_WritebackController_l84_132 = ((io_valuWrites_4_valid && io_vloadWrites_2_valid) && (io_valuWrites_4_payload_addr == io_vloadWrites_2_payload_addr));
  assign when_WritebackController_l84_133 = ((io_valuWrites_4_valid && io_vloadWrites_3_valid) && (io_valuWrites_4_payload_addr == io_vloadWrites_3_payload_addr));
  assign when_WritebackController_l84_134 = ((io_valuWrites_4_valid && io_vloadWrites_4_valid) && (io_valuWrites_4_payload_addr == io_vloadWrites_4_payload_addr));
  assign when_WritebackController_l84_135 = ((io_valuWrites_4_valid && io_vloadWrites_5_valid) && (io_valuWrites_4_payload_addr == io_vloadWrites_5_payload_addr));
  assign when_WritebackController_l84_136 = ((io_valuWrites_4_valid && io_vloadWrites_6_valid) && (io_valuWrites_4_payload_addr == io_vloadWrites_6_payload_addr));
  assign when_WritebackController_l84_137 = ((io_valuWrites_4_valid && io_vloadWrites_7_valid) && (io_valuWrites_4_payload_addr == io_vloadWrites_7_payload_addr));
  assign when_WritebackController_l84_138 = ((io_valuWrites_4_valid && io_flowScalarWrite_valid) && (io_valuWrites_4_payload_addr == io_flowScalarWrite_payload_addr));
  assign when_WritebackController_l84_139 = ((io_valuWrites_4_valid && io_flowVectorWrites_0_valid) && (io_valuWrites_4_payload_addr == io_flowVectorWrites_0_payload_addr));
  assign when_WritebackController_l84_140 = ((io_valuWrites_4_valid && io_flowVectorWrites_1_valid) && (io_valuWrites_4_payload_addr == io_flowVectorWrites_1_payload_addr));
  assign when_WritebackController_l84_141 = ((io_valuWrites_4_valid && io_flowVectorWrites_2_valid) && (io_valuWrites_4_payload_addr == io_flowVectorWrites_2_payload_addr));
  assign when_WritebackController_l84_142 = ((io_valuWrites_4_valid && io_flowVectorWrites_3_valid) && (io_valuWrites_4_payload_addr == io_flowVectorWrites_3_payload_addr));
  assign when_WritebackController_l84_143 = ((io_valuWrites_4_valid && io_flowVectorWrites_4_valid) && (io_valuWrites_4_payload_addr == io_flowVectorWrites_4_payload_addr));
  assign when_WritebackController_l84_144 = ((io_valuWrites_4_valid && io_flowVectorWrites_5_valid) && (io_valuWrites_4_payload_addr == io_flowVectorWrites_5_payload_addr));
  assign when_WritebackController_l84_145 = ((io_valuWrites_4_valid && io_flowVectorWrites_6_valid) && (io_valuWrites_4_payload_addr == io_flowVectorWrites_6_payload_addr));
  assign when_WritebackController_l84_146 = ((io_valuWrites_4_valid && io_flowVectorWrites_7_valid) && (io_valuWrites_4_payload_addr == io_flowVectorWrites_7_payload_addr));
  assign when_WritebackController_l84_147 = ((io_valuWrites_5_valid && io_valuWrites_6_valid) && (io_valuWrites_5_payload_addr == io_valuWrites_6_payload_addr));
  assign when_WritebackController_l84_148 = ((io_valuWrites_5_valid && io_valuWrites_7_valid) && (io_valuWrites_5_payload_addr == io_valuWrites_7_payload_addr));
  assign when_WritebackController_l84_149 = ((io_valuWrites_5_valid && io_loadWrites_0_valid) && (io_valuWrites_5_payload_addr == io_loadWrites_0_payload_addr));
  assign when_WritebackController_l84_150 = ((io_valuWrites_5_valid && io_constWrites_0_valid) && (io_valuWrites_5_payload_addr == io_constWrites_0_payload_addr));
  assign when_WritebackController_l84_151 = ((io_valuWrites_5_valid && io_vloadWrites_0_valid) && (io_valuWrites_5_payload_addr == io_vloadWrites_0_payload_addr));
  assign when_WritebackController_l84_152 = ((io_valuWrites_5_valid && io_vloadWrites_1_valid) && (io_valuWrites_5_payload_addr == io_vloadWrites_1_payload_addr));
  assign when_WritebackController_l84_153 = ((io_valuWrites_5_valid && io_vloadWrites_2_valid) && (io_valuWrites_5_payload_addr == io_vloadWrites_2_payload_addr));
  assign when_WritebackController_l84_154 = ((io_valuWrites_5_valid && io_vloadWrites_3_valid) && (io_valuWrites_5_payload_addr == io_vloadWrites_3_payload_addr));
  assign when_WritebackController_l84_155 = ((io_valuWrites_5_valid && io_vloadWrites_4_valid) && (io_valuWrites_5_payload_addr == io_vloadWrites_4_payload_addr));
  assign when_WritebackController_l84_156 = ((io_valuWrites_5_valid && io_vloadWrites_5_valid) && (io_valuWrites_5_payload_addr == io_vloadWrites_5_payload_addr));
  assign when_WritebackController_l84_157 = ((io_valuWrites_5_valid && io_vloadWrites_6_valid) && (io_valuWrites_5_payload_addr == io_vloadWrites_6_payload_addr));
  assign when_WritebackController_l84_158 = ((io_valuWrites_5_valid && io_vloadWrites_7_valid) && (io_valuWrites_5_payload_addr == io_vloadWrites_7_payload_addr));
  assign when_WritebackController_l84_159 = ((io_valuWrites_5_valid && io_flowScalarWrite_valid) && (io_valuWrites_5_payload_addr == io_flowScalarWrite_payload_addr));
  assign when_WritebackController_l84_160 = ((io_valuWrites_5_valid && io_flowVectorWrites_0_valid) && (io_valuWrites_5_payload_addr == io_flowVectorWrites_0_payload_addr));
  assign when_WritebackController_l84_161 = ((io_valuWrites_5_valid && io_flowVectorWrites_1_valid) && (io_valuWrites_5_payload_addr == io_flowVectorWrites_1_payload_addr));
  assign when_WritebackController_l84_162 = ((io_valuWrites_5_valid && io_flowVectorWrites_2_valid) && (io_valuWrites_5_payload_addr == io_flowVectorWrites_2_payload_addr));
  assign when_WritebackController_l84_163 = ((io_valuWrites_5_valid && io_flowVectorWrites_3_valid) && (io_valuWrites_5_payload_addr == io_flowVectorWrites_3_payload_addr));
  assign when_WritebackController_l84_164 = ((io_valuWrites_5_valid && io_flowVectorWrites_4_valid) && (io_valuWrites_5_payload_addr == io_flowVectorWrites_4_payload_addr));
  assign when_WritebackController_l84_165 = ((io_valuWrites_5_valid && io_flowVectorWrites_5_valid) && (io_valuWrites_5_payload_addr == io_flowVectorWrites_5_payload_addr));
  assign when_WritebackController_l84_166 = ((io_valuWrites_5_valid && io_flowVectorWrites_6_valid) && (io_valuWrites_5_payload_addr == io_flowVectorWrites_6_payload_addr));
  assign when_WritebackController_l84_167 = ((io_valuWrites_5_valid && io_flowVectorWrites_7_valid) && (io_valuWrites_5_payload_addr == io_flowVectorWrites_7_payload_addr));
  assign when_WritebackController_l84_168 = ((io_valuWrites_6_valid && io_valuWrites_7_valid) && (io_valuWrites_6_payload_addr == io_valuWrites_7_payload_addr));
  assign when_WritebackController_l84_169 = ((io_valuWrites_6_valid && io_loadWrites_0_valid) && (io_valuWrites_6_payload_addr == io_loadWrites_0_payload_addr));
  assign when_WritebackController_l84_170 = ((io_valuWrites_6_valid && io_constWrites_0_valid) && (io_valuWrites_6_payload_addr == io_constWrites_0_payload_addr));
  assign when_WritebackController_l84_171 = ((io_valuWrites_6_valid && io_vloadWrites_0_valid) && (io_valuWrites_6_payload_addr == io_vloadWrites_0_payload_addr));
  assign when_WritebackController_l84_172 = ((io_valuWrites_6_valid && io_vloadWrites_1_valid) && (io_valuWrites_6_payload_addr == io_vloadWrites_1_payload_addr));
  assign when_WritebackController_l84_173 = ((io_valuWrites_6_valid && io_vloadWrites_2_valid) && (io_valuWrites_6_payload_addr == io_vloadWrites_2_payload_addr));
  assign when_WritebackController_l84_174 = ((io_valuWrites_6_valid && io_vloadWrites_3_valid) && (io_valuWrites_6_payload_addr == io_vloadWrites_3_payload_addr));
  assign when_WritebackController_l84_175 = ((io_valuWrites_6_valid && io_vloadWrites_4_valid) && (io_valuWrites_6_payload_addr == io_vloadWrites_4_payload_addr));
  assign when_WritebackController_l84_176 = ((io_valuWrites_6_valid && io_vloadWrites_5_valid) && (io_valuWrites_6_payload_addr == io_vloadWrites_5_payload_addr));
  assign when_WritebackController_l84_177 = ((io_valuWrites_6_valid && io_vloadWrites_6_valid) && (io_valuWrites_6_payload_addr == io_vloadWrites_6_payload_addr));
  assign when_WritebackController_l84_178 = ((io_valuWrites_6_valid && io_vloadWrites_7_valid) && (io_valuWrites_6_payload_addr == io_vloadWrites_7_payload_addr));
  assign when_WritebackController_l84_179 = ((io_valuWrites_6_valid && io_flowScalarWrite_valid) && (io_valuWrites_6_payload_addr == io_flowScalarWrite_payload_addr));
  assign when_WritebackController_l84_180 = ((io_valuWrites_6_valid && io_flowVectorWrites_0_valid) && (io_valuWrites_6_payload_addr == io_flowVectorWrites_0_payload_addr));
  assign when_WritebackController_l84_181 = ((io_valuWrites_6_valid && io_flowVectorWrites_1_valid) && (io_valuWrites_6_payload_addr == io_flowVectorWrites_1_payload_addr));
  assign when_WritebackController_l84_182 = ((io_valuWrites_6_valid && io_flowVectorWrites_2_valid) && (io_valuWrites_6_payload_addr == io_flowVectorWrites_2_payload_addr));
  assign when_WritebackController_l84_183 = ((io_valuWrites_6_valid && io_flowVectorWrites_3_valid) && (io_valuWrites_6_payload_addr == io_flowVectorWrites_3_payload_addr));
  assign when_WritebackController_l84_184 = ((io_valuWrites_6_valid && io_flowVectorWrites_4_valid) && (io_valuWrites_6_payload_addr == io_flowVectorWrites_4_payload_addr));
  assign when_WritebackController_l84_185 = ((io_valuWrites_6_valid && io_flowVectorWrites_5_valid) && (io_valuWrites_6_payload_addr == io_flowVectorWrites_5_payload_addr));
  assign when_WritebackController_l84_186 = ((io_valuWrites_6_valid && io_flowVectorWrites_6_valid) && (io_valuWrites_6_payload_addr == io_flowVectorWrites_6_payload_addr));
  assign when_WritebackController_l84_187 = ((io_valuWrites_6_valid && io_flowVectorWrites_7_valid) && (io_valuWrites_6_payload_addr == io_flowVectorWrites_7_payload_addr));
  assign when_WritebackController_l84_188 = ((io_valuWrites_7_valid && io_loadWrites_0_valid) && (io_valuWrites_7_payload_addr == io_loadWrites_0_payload_addr));
  assign when_WritebackController_l84_189 = ((io_valuWrites_7_valid && io_constWrites_0_valid) && (io_valuWrites_7_payload_addr == io_constWrites_0_payload_addr));
  assign when_WritebackController_l84_190 = ((io_valuWrites_7_valid && io_vloadWrites_0_valid) && (io_valuWrites_7_payload_addr == io_vloadWrites_0_payload_addr));
  assign when_WritebackController_l84_191 = ((io_valuWrites_7_valid && io_vloadWrites_1_valid) && (io_valuWrites_7_payload_addr == io_vloadWrites_1_payload_addr));
  assign when_WritebackController_l84_192 = ((io_valuWrites_7_valid && io_vloadWrites_2_valid) && (io_valuWrites_7_payload_addr == io_vloadWrites_2_payload_addr));
  assign when_WritebackController_l84_193 = ((io_valuWrites_7_valid && io_vloadWrites_3_valid) && (io_valuWrites_7_payload_addr == io_vloadWrites_3_payload_addr));
  assign when_WritebackController_l84_194 = ((io_valuWrites_7_valid && io_vloadWrites_4_valid) && (io_valuWrites_7_payload_addr == io_vloadWrites_4_payload_addr));
  assign when_WritebackController_l84_195 = ((io_valuWrites_7_valid && io_vloadWrites_5_valid) && (io_valuWrites_7_payload_addr == io_vloadWrites_5_payload_addr));
  assign when_WritebackController_l84_196 = ((io_valuWrites_7_valid && io_vloadWrites_6_valid) && (io_valuWrites_7_payload_addr == io_vloadWrites_6_payload_addr));
  assign when_WritebackController_l84_197 = ((io_valuWrites_7_valid && io_vloadWrites_7_valid) && (io_valuWrites_7_payload_addr == io_vloadWrites_7_payload_addr));
  assign when_WritebackController_l84_198 = ((io_valuWrites_7_valid && io_flowScalarWrite_valid) && (io_valuWrites_7_payload_addr == io_flowScalarWrite_payload_addr));
  assign when_WritebackController_l84_199 = ((io_valuWrites_7_valid && io_flowVectorWrites_0_valid) && (io_valuWrites_7_payload_addr == io_flowVectorWrites_0_payload_addr));
  assign when_WritebackController_l84_200 = ((io_valuWrites_7_valid && io_flowVectorWrites_1_valid) && (io_valuWrites_7_payload_addr == io_flowVectorWrites_1_payload_addr));
  assign when_WritebackController_l84_201 = ((io_valuWrites_7_valid && io_flowVectorWrites_2_valid) && (io_valuWrites_7_payload_addr == io_flowVectorWrites_2_payload_addr));
  assign when_WritebackController_l84_202 = ((io_valuWrites_7_valid && io_flowVectorWrites_3_valid) && (io_valuWrites_7_payload_addr == io_flowVectorWrites_3_payload_addr));
  assign when_WritebackController_l84_203 = ((io_valuWrites_7_valid && io_flowVectorWrites_4_valid) && (io_valuWrites_7_payload_addr == io_flowVectorWrites_4_payload_addr));
  assign when_WritebackController_l84_204 = ((io_valuWrites_7_valid && io_flowVectorWrites_5_valid) && (io_valuWrites_7_payload_addr == io_flowVectorWrites_5_payload_addr));
  assign when_WritebackController_l84_205 = ((io_valuWrites_7_valid && io_flowVectorWrites_6_valid) && (io_valuWrites_7_payload_addr == io_flowVectorWrites_6_payload_addr));
  assign when_WritebackController_l84_206 = ((io_valuWrites_7_valid && io_flowVectorWrites_7_valid) && (io_valuWrites_7_payload_addr == io_flowVectorWrites_7_payload_addr));
  assign when_WritebackController_l84_207 = ((io_loadWrites_0_valid && io_constWrites_0_valid) && (io_loadWrites_0_payload_addr == io_constWrites_0_payload_addr));
  assign when_WritebackController_l84_208 = ((io_loadWrites_0_valid && io_vloadWrites_0_valid) && (io_loadWrites_0_payload_addr == io_vloadWrites_0_payload_addr));
  assign when_WritebackController_l84_209 = ((io_loadWrites_0_valid && io_vloadWrites_1_valid) && (io_loadWrites_0_payload_addr == io_vloadWrites_1_payload_addr));
  assign when_WritebackController_l84_210 = ((io_loadWrites_0_valid && io_vloadWrites_2_valid) && (io_loadWrites_0_payload_addr == io_vloadWrites_2_payload_addr));
  assign when_WritebackController_l84_211 = ((io_loadWrites_0_valid && io_vloadWrites_3_valid) && (io_loadWrites_0_payload_addr == io_vloadWrites_3_payload_addr));
  assign when_WritebackController_l84_212 = ((io_loadWrites_0_valid && io_vloadWrites_4_valid) && (io_loadWrites_0_payload_addr == io_vloadWrites_4_payload_addr));
  assign when_WritebackController_l84_213 = ((io_loadWrites_0_valid && io_vloadWrites_5_valid) && (io_loadWrites_0_payload_addr == io_vloadWrites_5_payload_addr));
  assign when_WritebackController_l84_214 = ((io_loadWrites_0_valid && io_vloadWrites_6_valid) && (io_loadWrites_0_payload_addr == io_vloadWrites_6_payload_addr));
  assign when_WritebackController_l84_215 = ((io_loadWrites_0_valid && io_vloadWrites_7_valid) && (io_loadWrites_0_payload_addr == io_vloadWrites_7_payload_addr));
  assign when_WritebackController_l84_216 = ((io_loadWrites_0_valid && io_flowScalarWrite_valid) && (io_loadWrites_0_payload_addr == io_flowScalarWrite_payload_addr));
  assign when_WritebackController_l84_217 = ((io_loadWrites_0_valid && io_flowVectorWrites_0_valid) && (io_loadWrites_0_payload_addr == io_flowVectorWrites_0_payload_addr));
  assign when_WritebackController_l84_218 = ((io_loadWrites_0_valid && io_flowVectorWrites_1_valid) && (io_loadWrites_0_payload_addr == io_flowVectorWrites_1_payload_addr));
  assign when_WritebackController_l84_219 = ((io_loadWrites_0_valid && io_flowVectorWrites_2_valid) && (io_loadWrites_0_payload_addr == io_flowVectorWrites_2_payload_addr));
  assign when_WritebackController_l84_220 = ((io_loadWrites_0_valid && io_flowVectorWrites_3_valid) && (io_loadWrites_0_payload_addr == io_flowVectorWrites_3_payload_addr));
  assign when_WritebackController_l84_221 = ((io_loadWrites_0_valid && io_flowVectorWrites_4_valid) && (io_loadWrites_0_payload_addr == io_flowVectorWrites_4_payload_addr));
  assign when_WritebackController_l84_222 = ((io_loadWrites_0_valid && io_flowVectorWrites_5_valid) && (io_loadWrites_0_payload_addr == io_flowVectorWrites_5_payload_addr));
  assign when_WritebackController_l84_223 = ((io_loadWrites_0_valid && io_flowVectorWrites_6_valid) && (io_loadWrites_0_payload_addr == io_flowVectorWrites_6_payload_addr));
  assign when_WritebackController_l84_224 = ((io_loadWrites_0_valid && io_flowVectorWrites_7_valid) && (io_loadWrites_0_payload_addr == io_flowVectorWrites_7_payload_addr));
  assign when_WritebackController_l84_225 = ((io_constWrites_0_valid && io_vloadWrites_0_valid) && (io_constWrites_0_payload_addr == io_vloadWrites_0_payload_addr));
  assign when_WritebackController_l84_226 = ((io_constWrites_0_valid && io_vloadWrites_1_valid) && (io_constWrites_0_payload_addr == io_vloadWrites_1_payload_addr));
  assign when_WritebackController_l84_227 = ((io_constWrites_0_valid && io_vloadWrites_2_valid) && (io_constWrites_0_payload_addr == io_vloadWrites_2_payload_addr));
  assign when_WritebackController_l84_228 = ((io_constWrites_0_valid && io_vloadWrites_3_valid) && (io_constWrites_0_payload_addr == io_vloadWrites_3_payload_addr));
  assign when_WritebackController_l84_229 = ((io_constWrites_0_valid && io_vloadWrites_4_valid) && (io_constWrites_0_payload_addr == io_vloadWrites_4_payload_addr));
  assign when_WritebackController_l84_230 = ((io_constWrites_0_valid && io_vloadWrites_5_valid) && (io_constWrites_0_payload_addr == io_vloadWrites_5_payload_addr));
  assign when_WritebackController_l84_231 = ((io_constWrites_0_valid && io_vloadWrites_6_valid) && (io_constWrites_0_payload_addr == io_vloadWrites_6_payload_addr));
  assign when_WritebackController_l84_232 = ((io_constWrites_0_valid && io_vloadWrites_7_valid) && (io_constWrites_0_payload_addr == io_vloadWrites_7_payload_addr));
  assign when_WritebackController_l84_233 = ((io_constWrites_0_valid && io_flowScalarWrite_valid) && (io_constWrites_0_payload_addr == io_flowScalarWrite_payload_addr));
  assign when_WritebackController_l84_234 = ((io_constWrites_0_valid && io_flowVectorWrites_0_valid) && (io_constWrites_0_payload_addr == io_flowVectorWrites_0_payload_addr));
  assign when_WritebackController_l84_235 = ((io_constWrites_0_valid && io_flowVectorWrites_1_valid) && (io_constWrites_0_payload_addr == io_flowVectorWrites_1_payload_addr));
  assign when_WritebackController_l84_236 = ((io_constWrites_0_valid && io_flowVectorWrites_2_valid) && (io_constWrites_0_payload_addr == io_flowVectorWrites_2_payload_addr));
  assign when_WritebackController_l84_237 = ((io_constWrites_0_valid && io_flowVectorWrites_3_valid) && (io_constWrites_0_payload_addr == io_flowVectorWrites_3_payload_addr));
  assign when_WritebackController_l84_238 = ((io_constWrites_0_valid && io_flowVectorWrites_4_valid) && (io_constWrites_0_payload_addr == io_flowVectorWrites_4_payload_addr));
  assign when_WritebackController_l84_239 = ((io_constWrites_0_valid && io_flowVectorWrites_5_valid) && (io_constWrites_0_payload_addr == io_flowVectorWrites_5_payload_addr));
  assign when_WritebackController_l84_240 = ((io_constWrites_0_valid && io_flowVectorWrites_6_valid) && (io_constWrites_0_payload_addr == io_flowVectorWrites_6_payload_addr));
  assign when_WritebackController_l84_241 = ((io_constWrites_0_valid && io_flowVectorWrites_7_valid) && (io_constWrites_0_payload_addr == io_flowVectorWrites_7_payload_addr));
  assign when_WritebackController_l84_242 = ((io_vloadWrites_0_valid && io_vloadWrites_1_valid) && (io_vloadWrites_0_payload_addr == io_vloadWrites_1_payload_addr));
  assign when_WritebackController_l84_243 = ((io_vloadWrites_0_valid && io_vloadWrites_2_valid) && (io_vloadWrites_0_payload_addr == io_vloadWrites_2_payload_addr));
  assign when_WritebackController_l84_244 = ((io_vloadWrites_0_valid && io_vloadWrites_3_valid) && (io_vloadWrites_0_payload_addr == io_vloadWrites_3_payload_addr));
  assign when_WritebackController_l84_245 = ((io_vloadWrites_0_valid && io_vloadWrites_4_valid) && (io_vloadWrites_0_payload_addr == io_vloadWrites_4_payload_addr));
  assign when_WritebackController_l84_246 = ((io_vloadWrites_0_valid && io_vloadWrites_5_valid) && (io_vloadWrites_0_payload_addr == io_vloadWrites_5_payload_addr));
  assign when_WritebackController_l84_247 = ((io_vloadWrites_0_valid && io_vloadWrites_6_valid) && (io_vloadWrites_0_payload_addr == io_vloadWrites_6_payload_addr));
  assign when_WritebackController_l84_248 = ((io_vloadWrites_0_valid && io_vloadWrites_7_valid) && (io_vloadWrites_0_payload_addr == io_vloadWrites_7_payload_addr));
  assign when_WritebackController_l84_249 = ((io_vloadWrites_0_valid && io_flowScalarWrite_valid) && (io_vloadWrites_0_payload_addr == io_flowScalarWrite_payload_addr));
  assign when_WritebackController_l84_250 = ((io_vloadWrites_0_valid && io_flowVectorWrites_0_valid) && (io_vloadWrites_0_payload_addr == io_flowVectorWrites_0_payload_addr));
  assign when_WritebackController_l84_251 = ((io_vloadWrites_0_valid && io_flowVectorWrites_1_valid) && (io_vloadWrites_0_payload_addr == io_flowVectorWrites_1_payload_addr));
  assign when_WritebackController_l84_252 = ((io_vloadWrites_0_valid && io_flowVectorWrites_2_valid) && (io_vloadWrites_0_payload_addr == io_flowVectorWrites_2_payload_addr));
  assign when_WritebackController_l84_253 = ((io_vloadWrites_0_valid && io_flowVectorWrites_3_valid) && (io_vloadWrites_0_payload_addr == io_flowVectorWrites_3_payload_addr));
  assign when_WritebackController_l84_254 = ((io_vloadWrites_0_valid && io_flowVectorWrites_4_valid) && (io_vloadWrites_0_payload_addr == io_flowVectorWrites_4_payload_addr));
  assign when_WritebackController_l84_255 = ((io_vloadWrites_0_valid && io_flowVectorWrites_5_valid) && (io_vloadWrites_0_payload_addr == io_flowVectorWrites_5_payload_addr));
  assign when_WritebackController_l84_256 = ((io_vloadWrites_0_valid && io_flowVectorWrites_6_valid) && (io_vloadWrites_0_payload_addr == io_flowVectorWrites_6_payload_addr));
  assign when_WritebackController_l84_257 = ((io_vloadWrites_0_valid && io_flowVectorWrites_7_valid) && (io_vloadWrites_0_payload_addr == io_flowVectorWrites_7_payload_addr));
  assign when_WritebackController_l84_258 = ((io_vloadWrites_1_valid && io_vloadWrites_2_valid) && (io_vloadWrites_1_payload_addr == io_vloadWrites_2_payload_addr));
  assign when_WritebackController_l84_259 = ((io_vloadWrites_1_valid && io_vloadWrites_3_valid) && (io_vloadWrites_1_payload_addr == io_vloadWrites_3_payload_addr));
  assign when_WritebackController_l84_260 = ((io_vloadWrites_1_valid && io_vloadWrites_4_valid) && (io_vloadWrites_1_payload_addr == io_vloadWrites_4_payload_addr));
  assign when_WritebackController_l84_261 = ((io_vloadWrites_1_valid && io_vloadWrites_5_valid) && (io_vloadWrites_1_payload_addr == io_vloadWrites_5_payload_addr));
  assign when_WritebackController_l84_262 = ((io_vloadWrites_1_valid && io_vloadWrites_6_valid) && (io_vloadWrites_1_payload_addr == io_vloadWrites_6_payload_addr));
  assign when_WritebackController_l84_263 = ((io_vloadWrites_1_valid && io_vloadWrites_7_valid) && (io_vloadWrites_1_payload_addr == io_vloadWrites_7_payload_addr));
  assign when_WritebackController_l84_264 = ((io_vloadWrites_1_valid && io_flowScalarWrite_valid) && (io_vloadWrites_1_payload_addr == io_flowScalarWrite_payload_addr));
  assign when_WritebackController_l84_265 = ((io_vloadWrites_1_valid && io_flowVectorWrites_0_valid) && (io_vloadWrites_1_payload_addr == io_flowVectorWrites_0_payload_addr));
  assign when_WritebackController_l84_266 = ((io_vloadWrites_1_valid && io_flowVectorWrites_1_valid) && (io_vloadWrites_1_payload_addr == io_flowVectorWrites_1_payload_addr));
  assign when_WritebackController_l84_267 = ((io_vloadWrites_1_valid && io_flowVectorWrites_2_valid) && (io_vloadWrites_1_payload_addr == io_flowVectorWrites_2_payload_addr));
  assign when_WritebackController_l84_268 = ((io_vloadWrites_1_valid && io_flowVectorWrites_3_valid) && (io_vloadWrites_1_payload_addr == io_flowVectorWrites_3_payload_addr));
  assign when_WritebackController_l84_269 = ((io_vloadWrites_1_valid && io_flowVectorWrites_4_valid) && (io_vloadWrites_1_payload_addr == io_flowVectorWrites_4_payload_addr));
  assign when_WritebackController_l84_270 = ((io_vloadWrites_1_valid && io_flowVectorWrites_5_valid) && (io_vloadWrites_1_payload_addr == io_flowVectorWrites_5_payload_addr));
  assign when_WritebackController_l84_271 = ((io_vloadWrites_1_valid && io_flowVectorWrites_6_valid) && (io_vloadWrites_1_payload_addr == io_flowVectorWrites_6_payload_addr));
  assign when_WritebackController_l84_272 = ((io_vloadWrites_1_valid && io_flowVectorWrites_7_valid) && (io_vloadWrites_1_payload_addr == io_flowVectorWrites_7_payload_addr));
  assign when_WritebackController_l84_273 = ((io_vloadWrites_2_valid && io_vloadWrites_3_valid) && (io_vloadWrites_2_payload_addr == io_vloadWrites_3_payload_addr));
  assign when_WritebackController_l84_274 = ((io_vloadWrites_2_valid && io_vloadWrites_4_valid) && (io_vloadWrites_2_payload_addr == io_vloadWrites_4_payload_addr));
  assign when_WritebackController_l84_275 = ((io_vloadWrites_2_valid && io_vloadWrites_5_valid) && (io_vloadWrites_2_payload_addr == io_vloadWrites_5_payload_addr));
  assign when_WritebackController_l84_276 = ((io_vloadWrites_2_valid && io_vloadWrites_6_valid) && (io_vloadWrites_2_payload_addr == io_vloadWrites_6_payload_addr));
  assign when_WritebackController_l84_277 = ((io_vloadWrites_2_valid && io_vloadWrites_7_valid) && (io_vloadWrites_2_payload_addr == io_vloadWrites_7_payload_addr));
  assign when_WritebackController_l84_278 = ((io_vloadWrites_2_valid && io_flowScalarWrite_valid) && (io_vloadWrites_2_payload_addr == io_flowScalarWrite_payload_addr));
  assign when_WritebackController_l84_279 = ((io_vloadWrites_2_valid && io_flowVectorWrites_0_valid) && (io_vloadWrites_2_payload_addr == io_flowVectorWrites_0_payload_addr));
  assign when_WritebackController_l84_280 = ((io_vloadWrites_2_valid && io_flowVectorWrites_1_valid) && (io_vloadWrites_2_payload_addr == io_flowVectorWrites_1_payload_addr));
  assign when_WritebackController_l84_281 = ((io_vloadWrites_2_valid && io_flowVectorWrites_2_valid) && (io_vloadWrites_2_payload_addr == io_flowVectorWrites_2_payload_addr));
  assign when_WritebackController_l84_282 = ((io_vloadWrites_2_valid && io_flowVectorWrites_3_valid) && (io_vloadWrites_2_payload_addr == io_flowVectorWrites_3_payload_addr));
  assign when_WritebackController_l84_283 = ((io_vloadWrites_2_valid && io_flowVectorWrites_4_valid) && (io_vloadWrites_2_payload_addr == io_flowVectorWrites_4_payload_addr));
  assign when_WritebackController_l84_284 = ((io_vloadWrites_2_valid && io_flowVectorWrites_5_valid) && (io_vloadWrites_2_payload_addr == io_flowVectorWrites_5_payload_addr));
  assign when_WritebackController_l84_285 = ((io_vloadWrites_2_valid && io_flowVectorWrites_6_valid) && (io_vloadWrites_2_payload_addr == io_flowVectorWrites_6_payload_addr));
  assign when_WritebackController_l84_286 = ((io_vloadWrites_2_valid && io_flowVectorWrites_7_valid) && (io_vloadWrites_2_payload_addr == io_flowVectorWrites_7_payload_addr));
  assign when_WritebackController_l84_287 = ((io_vloadWrites_3_valid && io_vloadWrites_4_valid) && (io_vloadWrites_3_payload_addr == io_vloadWrites_4_payload_addr));
  assign when_WritebackController_l84_288 = ((io_vloadWrites_3_valid && io_vloadWrites_5_valid) && (io_vloadWrites_3_payload_addr == io_vloadWrites_5_payload_addr));
  assign when_WritebackController_l84_289 = ((io_vloadWrites_3_valid && io_vloadWrites_6_valid) && (io_vloadWrites_3_payload_addr == io_vloadWrites_6_payload_addr));
  assign when_WritebackController_l84_290 = ((io_vloadWrites_3_valid && io_vloadWrites_7_valid) && (io_vloadWrites_3_payload_addr == io_vloadWrites_7_payload_addr));
  assign when_WritebackController_l84_291 = ((io_vloadWrites_3_valid && io_flowScalarWrite_valid) && (io_vloadWrites_3_payload_addr == io_flowScalarWrite_payload_addr));
  assign when_WritebackController_l84_292 = ((io_vloadWrites_3_valid && io_flowVectorWrites_0_valid) && (io_vloadWrites_3_payload_addr == io_flowVectorWrites_0_payload_addr));
  assign when_WritebackController_l84_293 = ((io_vloadWrites_3_valid && io_flowVectorWrites_1_valid) && (io_vloadWrites_3_payload_addr == io_flowVectorWrites_1_payload_addr));
  assign when_WritebackController_l84_294 = ((io_vloadWrites_3_valid && io_flowVectorWrites_2_valid) && (io_vloadWrites_3_payload_addr == io_flowVectorWrites_2_payload_addr));
  assign when_WritebackController_l84_295 = ((io_vloadWrites_3_valid && io_flowVectorWrites_3_valid) && (io_vloadWrites_3_payload_addr == io_flowVectorWrites_3_payload_addr));
  assign when_WritebackController_l84_296 = ((io_vloadWrites_3_valid && io_flowVectorWrites_4_valid) && (io_vloadWrites_3_payload_addr == io_flowVectorWrites_4_payload_addr));
  assign when_WritebackController_l84_297 = ((io_vloadWrites_3_valid && io_flowVectorWrites_5_valid) && (io_vloadWrites_3_payload_addr == io_flowVectorWrites_5_payload_addr));
  assign when_WritebackController_l84_298 = ((io_vloadWrites_3_valid && io_flowVectorWrites_6_valid) && (io_vloadWrites_3_payload_addr == io_flowVectorWrites_6_payload_addr));
  assign when_WritebackController_l84_299 = ((io_vloadWrites_3_valid && io_flowVectorWrites_7_valid) && (io_vloadWrites_3_payload_addr == io_flowVectorWrites_7_payload_addr));
  assign when_WritebackController_l84_300 = ((io_vloadWrites_4_valid && io_vloadWrites_5_valid) && (io_vloadWrites_4_payload_addr == io_vloadWrites_5_payload_addr));
  assign when_WritebackController_l84_301 = ((io_vloadWrites_4_valid && io_vloadWrites_6_valid) && (io_vloadWrites_4_payload_addr == io_vloadWrites_6_payload_addr));
  assign when_WritebackController_l84_302 = ((io_vloadWrites_4_valid && io_vloadWrites_7_valid) && (io_vloadWrites_4_payload_addr == io_vloadWrites_7_payload_addr));
  assign when_WritebackController_l84_303 = ((io_vloadWrites_4_valid && io_flowScalarWrite_valid) && (io_vloadWrites_4_payload_addr == io_flowScalarWrite_payload_addr));
  assign when_WritebackController_l84_304 = ((io_vloadWrites_4_valid && io_flowVectorWrites_0_valid) && (io_vloadWrites_4_payload_addr == io_flowVectorWrites_0_payload_addr));
  assign when_WritebackController_l84_305 = ((io_vloadWrites_4_valid && io_flowVectorWrites_1_valid) && (io_vloadWrites_4_payload_addr == io_flowVectorWrites_1_payload_addr));
  assign when_WritebackController_l84_306 = ((io_vloadWrites_4_valid && io_flowVectorWrites_2_valid) && (io_vloadWrites_4_payload_addr == io_flowVectorWrites_2_payload_addr));
  assign when_WritebackController_l84_307 = ((io_vloadWrites_4_valid && io_flowVectorWrites_3_valid) && (io_vloadWrites_4_payload_addr == io_flowVectorWrites_3_payload_addr));
  assign when_WritebackController_l84_308 = ((io_vloadWrites_4_valid && io_flowVectorWrites_4_valid) && (io_vloadWrites_4_payload_addr == io_flowVectorWrites_4_payload_addr));
  assign when_WritebackController_l84_309 = ((io_vloadWrites_4_valid && io_flowVectorWrites_5_valid) && (io_vloadWrites_4_payload_addr == io_flowVectorWrites_5_payload_addr));
  assign when_WritebackController_l84_310 = ((io_vloadWrites_4_valid && io_flowVectorWrites_6_valid) && (io_vloadWrites_4_payload_addr == io_flowVectorWrites_6_payload_addr));
  assign when_WritebackController_l84_311 = ((io_vloadWrites_4_valid && io_flowVectorWrites_7_valid) && (io_vloadWrites_4_payload_addr == io_flowVectorWrites_7_payload_addr));
  assign when_WritebackController_l84_312 = ((io_vloadWrites_5_valid && io_vloadWrites_6_valid) && (io_vloadWrites_5_payload_addr == io_vloadWrites_6_payload_addr));
  assign when_WritebackController_l84_313 = ((io_vloadWrites_5_valid && io_vloadWrites_7_valid) && (io_vloadWrites_5_payload_addr == io_vloadWrites_7_payload_addr));
  assign when_WritebackController_l84_314 = ((io_vloadWrites_5_valid && io_flowScalarWrite_valid) && (io_vloadWrites_5_payload_addr == io_flowScalarWrite_payload_addr));
  assign when_WritebackController_l84_315 = ((io_vloadWrites_5_valid && io_flowVectorWrites_0_valid) && (io_vloadWrites_5_payload_addr == io_flowVectorWrites_0_payload_addr));
  assign when_WritebackController_l84_316 = ((io_vloadWrites_5_valid && io_flowVectorWrites_1_valid) && (io_vloadWrites_5_payload_addr == io_flowVectorWrites_1_payload_addr));
  assign when_WritebackController_l84_317 = ((io_vloadWrites_5_valid && io_flowVectorWrites_2_valid) && (io_vloadWrites_5_payload_addr == io_flowVectorWrites_2_payload_addr));
  assign when_WritebackController_l84_318 = ((io_vloadWrites_5_valid && io_flowVectorWrites_3_valid) && (io_vloadWrites_5_payload_addr == io_flowVectorWrites_3_payload_addr));
  assign when_WritebackController_l84_319 = ((io_vloadWrites_5_valid && io_flowVectorWrites_4_valid) && (io_vloadWrites_5_payload_addr == io_flowVectorWrites_4_payload_addr));
  assign when_WritebackController_l84_320 = ((io_vloadWrites_5_valid && io_flowVectorWrites_5_valid) && (io_vloadWrites_5_payload_addr == io_flowVectorWrites_5_payload_addr));
  assign when_WritebackController_l84_321 = ((io_vloadWrites_5_valid && io_flowVectorWrites_6_valid) && (io_vloadWrites_5_payload_addr == io_flowVectorWrites_6_payload_addr));
  assign when_WritebackController_l84_322 = ((io_vloadWrites_5_valid && io_flowVectorWrites_7_valid) && (io_vloadWrites_5_payload_addr == io_flowVectorWrites_7_payload_addr));
  assign when_WritebackController_l84_323 = ((io_vloadWrites_6_valid && io_vloadWrites_7_valid) && (io_vloadWrites_6_payload_addr == io_vloadWrites_7_payload_addr));
  assign when_WritebackController_l84_324 = ((io_vloadWrites_6_valid && io_flowScalarWrite_valid) && (io_vloadWrites_6_payload_addr == io_flowScalarWrite_payload_addr));
  assign when_WritebackController_l84_325 = ((io_vloadWrites_6_valid && io_flowVectorWrites_0_valid) && (io_vloadWrites_6_payload_addr == io_flowVectorWrites_0_payload_addr));
  assign when_WritebackController_l84_326 = ((io_vloadWrites_6_valid && io_flowVectorWrites_1_valid) && (io_vloadWrites_6_payload_addr == io_flowVectorWrites_1_payload_addr));
  assign when_WritebackController_l84_327 = ((io_vloadWrites_6_valid && io_flowVectorWrites_2_valid) && (io_vloadWrites_6_payload_addr == io_flowVectorWrites_2_payload_addr));
  assign when_WritebackController_l84_328 = ((io_vloadWrites_6_valid && io_flowVectorWrites_3_valid) && (io_vloadWrites_6_payload_addr == io_flowVectorWrites_3_payload_addr));
  assign when_WritebackController_l84_329 = ((io_vloadWrites_6_valid && io_flowVectorWrites_4_valid) && (io_vloadWrites_6_payload_addr == io_flowVectorWrites_4_payload_addr));
  assign when_WritebackController_l84_330 = ((io_vloadWrites_6_valid && io_flowVectorWrites_5_valid) && (io_vloadWrites_6_payload_addr == io_flowVectorWrites_5_payload_addr));
  assign when_WritebackController_l84_331 = ((io_vloadWrites_6_valid && io_flowVectorWrites_6_valid) && (io_vloadWrites_6_payload_addr == io_flowVectorWrites_6_payload_addr));
  assign when_WritebackController_l84_332 = ((io_vloadWrites_6_valid && io_flowVectorWrites_7_valid) && (io_vloadWrites_6_payload_addr == io_flowVectorWrites_7_payload_addr));
  assign when_WritebackController_l84_333 = ((io_vloadWrites_7_valid && io_flowScalarWrite_valid) && (io_vloadWrites_7_payload_addr == io_flowScalarWrite_payload_addr));
  assign when_WritebackController_l84_334 = ((io_vloadWrites_7_valid && io_flowVectorWrites_0_valid) && (io_vloadWrites_7_payload_addr == io_flowVectorWrites_0_payload_addr));
  assign when_WritebackController_l84_335 = ((io_vloadWrites_7_valid && io_flowVectorWrites_1_valid) && (io_vloadWrites_7_payload_addr == io_flowVectorWrites_1_payload_addr));
  assign when_WritebackController_l84_336 = ((io_vloadWrites_7_valid && io_flowVectorWrites_2_valid) && (io_vloadWrites_7_payload_addr == io_flowVectorWrites_2_payload_addr));
  assign when_WritebackController_l84_337 = ((io_vloadWrites_7_valid && io_flowVectorWrites_3_valid) && (io_vloadWrites_7_payload_addr == io_flowVectorWrites_3_payload_addr));
  assign when_WritebackController_l84_338 = ((io_vloadWrites_7_valid && io_flowVectorWrites_4_valid) && (io_vloadWrites_7_payload_addr == io_flowVectorWrites_4_payload_addr));
  assign when_WritebackController_l84_339 = ((io_vloadWrites_7_valid && io_flowVectorWrites_5_valid) && (io_vloadWrites_7_payload_addr == io_flowVectorWrites_5_payload_addr));
  assign when_WritebackController_l84_340 = ((io_vloadWrites_7_valid && io_flowVectorWrites_6_valid) && (io_vloadWrites_7_payload_addr == io_flowVectorWrites_6_payload_addr));
  assign when_WritebackController_l84_341 = ((io_vloadWrites_7_valid && io_flowVectorWrites_7_valid) && (io_vloadWrites_7_payload_addr == io_flowVectorWrites_7_payload_addr));
  assign when_WritebackController_l84_342 = ((io_flowScalarWrite_valid && io_flowVectorWrites_0_valid) && (io_flowScalarWrite_payload_addr == io_flowVectorWrites_0_payload_addr));
  assign when_WritebackController_l84_343 = ((io_flowScalarWrite_valid && io_flowVectorWrites_1_valid) && (io_flowScalarWrite_payload_addr == io_flowVectorWrites_1_payload_addr));
  assign when_WritebackController_l84_344 = ((io_flowScalarWrite_valid && io_flowVectorWrites_2_valid) && (io_flowScalarWrite_payload_addr == io_flowVectorWrites_2_payload_addr));
  assign when_WritebackController_l84_345 = ((io_flowScalarWrite_valid && io_flowVectorWrites_3_valid) && (io_flowScalarWrite_payload_addr == io_flowVectorWrites_3_payload_addr));
  assign when_WritebackController_l84_346 = ((io_flowScalarWrite_valid && io_flowVectorWrites_4_valid) && (io_flowScalarWrite_payload_addr == io_flowVectorWrites_4_payload_addr));
  assign when_WritebackController_l84_347 = ((io_flowScalarWrite_valid && io_flowVectorWrites_5_valid) && (io_flowScalarWrite_payload_addr == io_flowVectorWrites_5_payload_addr));
  assign when_WritebackController_l84_348 = ((io_flowScalarWrite_valid && io_flowVectorWrites_6_valid) && (io_flowScalarWrite_payload_addr == io_flowVectorWrites_6_payload_addr));
  assign when_WritebackController_l84_349 = ((io_flowScalarWrite_valid && io_flowVectorWrites_7_valid) && (io_flowScalarWrite_payload_addr == io_flowVectorWrites_7_payload_addr));
  assign when_WritebackController_l84_350 = ((io_flowVectorWrites_0_valid && io_flowVectorWrites_1_valid) && (io_flowVectorWrites_0_payload_addr == io_flowVectorWrites_1_payload_addr));
  assign when_WritebackController_l84_351 = ((io_flowVectorWrites_0_valid && io_flowVectorWrites_2_valid) && (io_flowVectorWrites_0_payload_addr == io_flowVectorWrites_2_payload_addr));
  assign when_WritebackController_l84_352 = ((io_flowVectorWrites_0_valid && io_flowVectorWrites_3_valid) && (io_flowVectorWrites_0_payload_addr == io_flowVectorWrites_3_payload_addr));
  assign when_WritebackController_l84_353 = ((io_flowVectorWrites_0_valid && io_flowVectorWrites_4_valid) && (io_flowVectorWrites_0_payload_addr == io_flowVectorWrites_4_payload_addr));
  assign when_WritebackController_l84_354 = ((io_flowVectorWrites_0_valid && io_flowVectorWrites_5_valid) && (io_flowVectorWrites_0_payload_addr == io_flowVectorWrites_5_payload_addr));
  assign when_WritebackController_l84_355 = ((io_flowVectorWrites_0_valid && io_flowVectorWrites_6_valid) && (io_flowVectorWrites_0_payload_addr == io_flowVectorWrites_6_payload_addr));
  assign when_WritebackController_l84_356 = ((io_flowVectorWrites_0_valid && io_flowVectorWrites_7_valid) && (io_flowVectorWrites_0_payload_addr == io_flowVectorWrites_7_payload_addr));
  assign when_WritebackController_l84_357 = ((io_flowVectorWrites_1_valid && io_flowVectorWrites_2_valid) && (io_flowVectorWrites_1_payload_addr == io_flowVectorWrites_2_payload_addr));
  assign when_WritebackController_l84_358 = ((io_flowVectorWrites_1_valid && io_flowVectorWrites_3_valid) && (io_flowVectorWrites_1_payload_addr == io_flowVectorWrites_3_payload_addr));
  assign when_WritebackController_l84_359 = ((io_flowVectorWrites_1_valid && io_flowVectorWrites_4_valid) && (io_flowVectorWrites_1_payload_addr == io_flowVectorWrites_4_payload_addr));
  assign when_WritebackController_l84_360 = ((io_flowVectorWrites_1_valid && io_flowVectorWrites_5_valid) && (io_flowVectorWrites_1_payload_addr == io_flowVectorWrites_5_payload_addr));
  assign when_WritebackController_l84_361 = ((io_flowVectorWrites_1_valid && io_flowVectorWrites_6_valid) && (io_flowVectorWrites_1_payload_addr == io_flowVectorWrites_6_payload_addr));
  assign when_WritebackController_l84_362 = ((io_flowVectorWrites_1_valid && io_flowVectorWrites_7_valid) && (io_flowVectorWrites_1_payload_addr == io_flowVectorWrites_7_payload_addr));
  assign when_WritebackController_l84_363 = ((io_flowVectorWrites_2_valid && io_flowVectorWrites_3_valid) && (io_flowVectorWrites_2_payload_addr == io_flowVectorWrites_3_payload_addr));
  assign when_WritebackController_l84_364 = ((io_flowVectorWrites_2_valid && io_flowVectorWrites_4_valid) && (io_flowVectorWrites_2_payload_addr == io_flowVectorWrites_4_payload_addr));
  assign when_WritebackController_l84_365 = ((io_flowVectorWrites_2_valid && io_flowVectorWrites_5_valid) && (io_flowVectorWrites_2_payload_addr == io_flowVectorWrites_5_payload_addr));
  assign when_WritebackController_l84_366 = ((io_flowVectorWrites_2_valid && io_flowVectorWrites_6_valid) && (io_flowVectorWrites_2_payload_addr == io_flowVectorWrites_6_payload_addr));
  assign when_WritebackController_l84_367 = ((io_flowVectorWrites_2_valid && io_flowVectorWrites_7_valid) && (io_flowVectorWrites_2_payload_addr == io_flowVectorWrites_7_payload_addr));
  assign when_WritebackController_l84_368 = ((io_flowVectorWrites_3_valid && io_flowVectorWrites_4_valid) && (io_flowVectorWrites_3_payload_addr == io_flowVectorWrites_4_payload_addr));
  assign when_WritebackController_l84_369 = ((io_flowVectorWrites_3_valid && io_flowVectorWrites_5_valid) && (io_flowVectorWrites_3_payload_addr == io_flowVectorWrites_5_payload_addr));
  assign when_WritebackController_l84_370 = ((io_flowVectorWrites_3_valid && io_flowVectorWrites_6_valid) && (io_flowVectorWrites_3_payload_addr == io_flowVectorWrites_6_payload_addr));
  assign when_WritebackController_l84_371 = ((io_flowVectorWrites_3_valid && io_flowVectorWrites_7_valid) && (io_flowVectorWrites_3_payload_addr == io_flowVectorWrites_7_payload_addr));
  assign when_WritebackController_l84_372 = ((io_flowVectorWrites_4_valid && io_flowVectorWrites_5_valid) && (io_flowVectorWrites_4_payload_addr == io_flowVectorWrites_5_payload_addr));
  assign when_WritebackController_l84_373 = ((io_flowVectorWrites_4_valid && io_flowVectorWrites_6_valid) && (io_flowVectorWrites_4_payload_addr == io_flowVectorWrites_6_payload_addr));
  assign when_WritebackController_l84_374 = ((io_flowVectorWrites_4_valid && io_flowVectorWrites_7_valid) && (io_flowVectorWrites_4_payload_addr == io_flowVectorWrites_7_payload_addr));
  assign when_WritebackController_l84_375 = ((io_flowVectorWrites_5_valid && io_flowVectorWrites_6_valid) && (io_flowVectorWrites_5_payload_addr == io_flowVectorWrites_6_payload_addr));
  assign when_WritebackController_l84_376 = ((io_flowVectorWrites_5_valid && io_flowVectorWrites_7_valid) && (io_flowVectorWrites_5_payload_addr == io_flowVectorWrites_7_payload_addr));
  assign when_WritebackController_l84_377 = ((io_flowVectorWrites_6_valid && io_flowVectorWrites_7_valid) && (io_flowVectorWrites_6_payload_addr == io_flowVectorWrites_7_payload_addr));
  always @(posedge clk) begin
    if(reset) begin
    end else begin
      if(when_WritebackController_l84) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 0 and port 1 both writing to addr %x", io_aluWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_1) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 0 and port 2 both writing to addr %x", io_aluWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_2) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 0 and port 3 both writing to addr %x", io_aluWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_3) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 0 and port 4 both writing to addr %x", io_aluWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_4) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 0 and port 5 both writing to addr %x", io_aluWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_5) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 0 and port 6 both writing to addr %x", io_aluWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_6) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 0 and port 7 both writing to addr %x", io_aluWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_7) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 0 and port 8 both writing to addr %x", io_aluWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_8) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 0 and port 9 both writing to addr %x", io_aluWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_9) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 0 and port 10 both writing to addr %x", io_aluWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_10) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 0 and port 11 both writing to addr %x", io_aluWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_11) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 0 and port 12 both writing to addr %x", io_aluWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_12) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 0 and port 13 both writing to addr %x", io_aluWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_13) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 0 and port 14 both writing to addr %x", io_aluWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_14) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 0 and port 15 both writing to addr %x", io_aluWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_15) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 0 and port 16 both writing to addr %x", io_aluWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_16) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 0 and port 17 both writing to addr %x", io_aluWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_17) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 0 and port 18 both writing to addr %x", io_aluWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_18) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 0 and port 19 both writing to addr %x", io_aluWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_19) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 0 and port 20 both writing to addr %x", io_aluWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_20) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 0 and port 21 both writing to addr %x", io_aluWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_21) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 0 and port 22 both writing to addr %x", io_aluWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_22) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 0 and port 23 both writing to addr %x", io_aluWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_23) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 0 and port 24 both writing to addr %x", io_aluWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_24) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 0 and port 25 both writing to addr %x", io_aluWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_25) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 0 and port 26 both writing to addr %x", io_aluWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_26) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 0 and port 27 both writing to addr %x", io_aluWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_27) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 1 and port 2 both writing to addr %x", io_valuWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_28) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 1 and port 3 both writing to addr %x", io_valuWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_29) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 1 and port 4 both writing to addr %x", io_valuWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_30) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 1 and port 5 both writing to addr %x", io_valuWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_31) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 1 and port 6 both writing to addr %x", io_valuWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_32) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 1 and port 7 both writing to addr %x", io_valuWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_33) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 1 and port 8 both writing to addr %x", io_valuWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_34) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 1 and port 9 both writing to addr %x", io_valuWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_35) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 1 and port 10 both writing to addr %x", io_valuWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_36) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 1 and port 11 both writing to addr %x", io_valuWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_37) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 1 and port 12 both writing to addr %x", io_valuWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_38) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 1 and port 13 both writing to addr %x", io_valuWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_39) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 1 and port 14 both writing to addr %x", io_valuWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_40) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 1 and port 15 both writing to addr %x", io_valuWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_41) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 1 and port 16 both writing to addr %x", io_valuWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_42) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 1 and port 17 both writing to addr %x", io_valuWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_43) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 1 and port 18 both writing to addr %x", io_valuWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_44) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 1 and port 19 both writing to addr %x", io_valuWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_45) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 1 and port 20 both writing to addr %x", io_valuWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_46) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 1 and port 21 both writing to addr %x", io_valuWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_47) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 1 and port 22 both writing to addr %x", io_valuWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_48) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 1 and port 23 both writing to addr %x", io_valuWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_49) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 1 and port 24 both writing to addr %x", io_valuWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_50) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 1 and port 25 both writing to addr %x", io_valuWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_51) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 1 and port 26 both writing to addr %x", io_valuWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_52) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 1 and port 27 both writing to addr %x", io_valuWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_53) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 2 and port 3 both writing to addr %x", io_valuWrites_1_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_54) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 2 and port 4 both writing to addr %x", io_valuWrites_1_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_55) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 2 and port 5 both writing to addr %x", io_valuWrites_1_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_56) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 2 and port 6 both writing to addr %x", io_valuWrites_1_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_57) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 2 and port 7 both writing to addr %x", io_valuWrites_1_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_58) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 2 and port 8 both writing to addr %x", io_valuWrites_1_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_59) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 2 and port 9 both writing to addr %x", io_valuWrites_1_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_60) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 2 and port 10 both writing to addr %x", io_valuWrites_1_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_61) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 2 and port 11 both writing to addr %x", io_valuWrites_1_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_62) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 2 and port 12 both writing to addr %x", io_valuWrites_1_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_63) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 2 and port 13 both writing to addr %x", io_valuWrites_1_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_64) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 2 and port 14 both writing to addr %x", io_valuWrites_1_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_65) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 2 and port 15 both writing to addr %x", io_valuWrites_1_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_66) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 2 and port 16 both writing to addr %x", io_valuWrites_1_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_67) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 2 and port 17 both writing to addr %x", io_valuWrites_1_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_68) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 2 and port 18 both writing to addr %x", io_valuWrites_1_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_69) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 2 and port 19 both writing to addr %x", io_valuWrites_1_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_70) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 2 and port 20 both writing to addr %x", io_valuWrites_1_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_71) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 2 and port 21 both writing to addr %x", io_valuWrites_1_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_72) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 2 and port 22 both writing to addr %x", io_valuWrites_1_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_73) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 2 and port 23 both writing to addr %x", io_valuWrites_1_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_74) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 2 and port 24 both writing to addr %x", io_valuWrites_1_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_75) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 2 and port 25 both writing to addr %x", io_valuWrites_1_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_76) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 2 and port 26 both writing to addr %x", io_valuWrites_1_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_77) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 2 and port 27 both writing to addr %x", io_valuWrites_1_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_78) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 3 and port 4 both writing to addr %x", io_valuWrites_2_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_79) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 3 and port 5 both writing to addr %x", io_valuWrites_2_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_80) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 3 and port 6 both writing to addr %x", io_valuWrites_2_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_81) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 3 and port 7 both writing to addr %x", io_valuWrites_2_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_82) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 3 and port 8 both writing to addr %x", io_valuWrites_2_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_83) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 3 and port 9 both writing to addr %x", io_valuWrites_2_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_84) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 3 and port 10 both writing to addr %x", io_valuWrites_2_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_85) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 3 and port 11 both writing to addr %x", io_valuWrites_2_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_86) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 3 and port 12 both writing to addr %x", io_valuWrites_2_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_87) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 3 and port 13 both writing to addr %x", io_valuWrites_2_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_88) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 3 and port 14 both writing to addr %x", io_valuWrites_2_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_89) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 3 and port 15 both writing to addr %x", io_valuWrites_2_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_90) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 3 and port 16 both writing to addr %x", io_valuWrites_2_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_91) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 3 and port 17 both writing to addr %x", io_valuWrites_2_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_92) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 3 and port 18 both writing to addr %x", io_valuWrites_2_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_93) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 3 and port 19 both writing to addr %x", io_valuWrites_2_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_94) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 3 and port 20 both writing to addr %x", io_valuWrites_2_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_95) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 3 and port 21 both writing to addr %x", io_valuWrites_2_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_96) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 3 and port 22 both writing to addr %x", io_valuWrites_2_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_97) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 3 and port 23 both writing to addr %x", io_valuWrites_2_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_98) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 3 and port 24 both writing to addr %x", io_valuWrites_2_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_99) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 3 and port 25 both writing to addr %x", io_valuWrites_2_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_100) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 3 and port 26 both writing to addr %x", io_valuWrites_2_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_101) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 3 and port 27 both writing to addr %x", io_valuWrites_2_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_102) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 4 and port 5 both writing to addr %x", io_valuWrites_3_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_103) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 4 and port 6 both writing to addr %x", io_valuWrites_3_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_104) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 4 and port 7 both writing to addr %x", io_valuWrites_3_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_105) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 4 and port 8 both writing to addr %x", io_valuWrites_3_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_106) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 4 and port 9 both writing to addr %x", io_valuWrites_3_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_107) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 4 and port 10 both writing to addr %x", io_valuWrites_3_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_108) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 4 and port 11 both writing to addr %x", io_valuWrites_3_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_109) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 4 and port 12 both writing to addr %x", io_valuWrites_3_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_110) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 4 and port 13 both writing to addr %x", io_valuWrites_3_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_111) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 4 and port 14 both writing to addr %x", io_valuWrites_3_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_112) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 4 and port 15 both writing to addr %x", io_valuWrites_3_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_113) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 4 and port 16 both writing to addr %x", io_valuWrites_3_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_114) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 4 and port 17 both writing to addr %x", io_valuWrites_3_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_115) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 4 and port 18 both writing to addr %x", io_valuWrites_3_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_116) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 4 and port 19 both writing to addr %x", io_valuWrites_3_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_117) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 4 and port 20 both writing to addr %x", io_valuWrites_3_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_118) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 4 and port 21 both writing to addr %x", io_valuWrites_3_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_119) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 4 and port 22 both writing to addr %x", io_valuWrites_3_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_120) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 4 and port 23 both writing to addr %x", io_valuWrites_3_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_121) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 4 and port 24 both writing to addr %x", io_valuWrites_3_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_122) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 4 and port 25 both writing to addr %x", io_valuWrites_3_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_123) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 4 and port 26 both writing to addr %x", io_valuWrites_3_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_124) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 4 and port 27 both writing to addr %x", io_valuWrites_3_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_125) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 5 and port 6 both writing to addr %x", io_valuWrites_4_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_126) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 5 and port 7 both writing to addr %x", io_valuWrites_4_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_127) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 5 and port 8 both writing to addr %x", io_valuWrites_4_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_128) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 5 and port 9 both writing to addr %x", io_valuWrites_4_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_129) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 5 and port 10 both writing to addr %x", io_valuWrites_4_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_130) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 5 and port 11 both writing to addr %x", io_valuWrites_4_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_131) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 5 and port 12 both writing to addr %x", io_valuWrites_4_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_132) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 5 and port 13 both writing to addr %x", io_valuWrites_4_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_133) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 5 and port 14 both writing to addr %x", io_valuWrites_4_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_134) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 5 and port 15 both writing to addr %x", io_valuWrites_4_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_135) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 5 and port 16 both writing to addr %x", io_valuWrites_4_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_136) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 5 and port 17 both writing to addr %x", io_valuWrites_4_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_137) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 5 and port 18 both writing to addr %x", io_valuWrites_4_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_138) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 5 and port 19 both writing to addr %x", io_valuWrites_4_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_139) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 5 and port 20 both writing to addr %x", io_valuWrites_4_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_140) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 5 and port 21 both writing to addr %x", io_valuWrites_4_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_141) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 5 and port 22 both writing to addr %x", io_valuWrites_4_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_142) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 5 and port 23 both writing to addr %x", io_valuWrites_4_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_143) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 5 and port 24 both writing to addr %x", io_valuWrites_4_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_144) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 5 and port 25 both writing to addr %x", io_valuWrites_4_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_145) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 5 and port 26 both writing to addr %x", io_valuWrites_4_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_146) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 5 and port 27 both writing to addr %x", io_valuWrites_4_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_147) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 6 and port 7 both writing to addr %x", io_valuWrites_5_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_148) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 6 and port 8 both writing to addr %x", io_valuWrites_5_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_149) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 6 and port 9 both writing to addr %x", io_valuWrites_5_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_150) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 6 and port 10 both writing to addr %x", io_valuWrites_5_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_151) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 6 and port 11 both writing to addr %x", io_valuWrites_5_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_152) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 6 and port 12 both writing to addr %x", io_valuWrites_5_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_153) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 6 and port 13 both writing to addr %x", io_valuWrites_5_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_154) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 6 and port 14 both writing to addr %x", io_valuWrites_5_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_155) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 6 and port 15 both writing to addr %x", io_valuWrites_5_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_156) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 6 and port 16 both writing to addr %x", io_valuWrites_5_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_157) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 6 and port 17 both writing to addr %x", io_valuWrites_5_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_158) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 6 and port 18 both writing to addr %x", io_valuWrites_5_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_159) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 6 and port 19 both writing to addr %x", io_valuWrites_5_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_160) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 6 and port 20 both writing to addr %x", io_valuWrites_5_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_161) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 6 and port 21 both writing to addr %x", io_valuWrites_5_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_162) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 6 and port 22 both writing to addr %x", io_valuWrites_5_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_163) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 6 and port 23 both writing to addr %x", io_valuWrites_5_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_164) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 6 and port 24 both writing to addr %x", io_valuWrites_5_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_165) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 6 and port 25 both writing to addr %x", io_valuWrites_5_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_166) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 6 and port 26 both writing to addr %x", io_valuWrites_5_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_167) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 6 and port 27 both writing to addr %x", io_valuWrites_5_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_168) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 7 and port 8 both writing to addr %x", io_valuWrites_6_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_169) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 7 and port 9 both writing to addr %x", io_valuWrites_6_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_170) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 7 and port 10 both writing to addr %x", io_valuWrites_6_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_171) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 7 and port 11 both writing to addr %x", io_valuWrites_6_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_172) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 7 and port 12 both writing to addr %x", io_valuWrites_6_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_173) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 7 and port 13 both writing to addr %x", io_valuWrites_6_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_174) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 7 and port 14 both writing to addr %x", io_valuWrites_6_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_175) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 7 and port 15 both writing to addr %x", io_valuWrites_6_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_176) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 7 and port 16 both writing to addr %x", io_valuWrites_6_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_177) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 7 and port 17 both writing to addr %x", io_valuWrites_6_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_178) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 7 and port 18 both writing to addr %x", io_valuWrites_6_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_179) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 7 and port 19 both writing to addr %x", io_valuWrites_6_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_180) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 7 and port 20 both writing to addr %x", io_valuWrites_6_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_181) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 7 and port 21 both writing to addr %x", io_valuWrites_6_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_182) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 7 and port 22 both writing to addr %x", io_valuWrites_6_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_183) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 7 and port 23 both writing to addr %x", io_valuWrites_6_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_184) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 7 and port 24 both writing to addr %x", io_valuWrites_6_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_185) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 7 and port 25 both writing to addr %x", io_valuWrites_6_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_186) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 7 and port 26 both writing to addr %x", io_valuWrites_6_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_187) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 7 and port 27 both writing to addr %x", io_valuWrites_6_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_188) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 8 and port 9 both writing to addr %x", io_valuWrites_7_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_189) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 8 and port 10 both writing to addr %x", io_valuWrites_7_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_190) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 8 and port 11 both writing to addr %x", io_valuWrites_7_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_191) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 8 and port 12 both writing to addr %x", io_valuWrites_7_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_192) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 8 and port 13 both writing to addr %x", io_valuWrites_7_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_193) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 8 and port 14 both writing to addr %x", io_valuWrites_7_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_194) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 8 and port 15 both writing to addr %x", io_valuWrites_7_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_195) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 8 and port 16 both writing to addr %x", io_valuWrites_7_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_196) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 8 and port 17 both writing to addr %x", io_valuWrites_7_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_197) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 8 and port 18 both writing to addr %x", io_valuWrites_7_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_198) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 8 and port 19 both writing to addr %x", io_valuWrites_7_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_199) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 8 and port 20 both writing to addr %x", io_valuWrites_7_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_200) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 8 and port 21 both writing to addr %x", io_valuWrites_7_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_201) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 8 and port 22 both writing to addr %x", io_valuWrites_7_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_202) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 8 and port 23 both writing to addr %x", io_valuWrites_7_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_203) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 8 and port 24 both writing to addr %x", io_valuWrites_7_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_204) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 8 and port 25 both writing to addr %x", io_valuWrites_7_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_205) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 8 and port 26 both writing to addr %x", io_valuWrites_7_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_206) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 8 and port 27 both writing to addr %x", io_valuWrites_7_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_207) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 9 and port 10 both writing to addr %x", io_loadWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_208) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 9 and port 11 both writing to addr %x", io_loadWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_209) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 9 and port 12 both writing to addr %x", io_loadWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_210) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 9 and port 13 both writing to addr %x", io_loadWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_211) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 9 and port 14 both writing to addr %x", io_loadWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_212) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 9 and port 15 both writing to addr %x", io_loadWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_213) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 9 and port 16 both writing to addr %x", io_loadWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_214) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 9 and port 17 both writing to addr %x", io_loadWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_215) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 9 and port 18 both writing to addr %x", io_loadWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_216) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 9 and port 19 both writing to addr %x", io_loadWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_217) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 9 and port 20 both writing to addr %x", io_loadWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_218) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 9 and port 21 both writing to addr %x", io_loadWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_219) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 9 and port 22 both writing to addr %x", io_loadWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_220) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 9 and port 23 both writing to addr %x", io_loadWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_221) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 9 and port 24 both writing to addr %x", io_loadWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_222) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 9 and port 25 both writing to addr %x", io_loadWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_223) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 9 and port 26 both writing to addr %x", io_loadWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_224) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 9 and port 27 both writing to addr %x", io_loadWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_225) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 10 and port 11 both writing to addr %x", io_constWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_226) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 10 and port 12 both writing to addr %x", io_constWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_227) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 10 and port 13 both writing to addr %x", io_constWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_228) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 10 and port 14 both writing to addr %x", io_constWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_229) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 10 and port 15 both writing to addr %x", io_constWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_230) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 10 and port 16 both writing to addr %x", io_constWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_231) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 10 and port 17 both writing to addr %x", io_constWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_232) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 10 and port 18 both writing to addr %x", io_constWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_233) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 10 and port 19 both writing to addr %x", io_constWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_234) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 10 and port 20 both writing to addr %x", io_constWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_235) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 10 and port 21 both writing to addr %x", io_constWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_236) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 10 and port 22 both writing to addr %x", io_constWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_237) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 10 and port 23 both writing to addr %x", io_constWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_238) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 10 and port 24 both writing to addr %x", io_constWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_239) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 10 and port 25 both writing to addr %x", io_constWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_240) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 10 and port 26 both writing to addr %x", io_constWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_241) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 10 and port 27 both writing to addr %x", io_constWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_242) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 11 and port 12 both writing to addr %x", io_vloadWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_243) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 11 and port 13 both writing to addr %x", io_vloadWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_244) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 11 and port 14 both writing to addr %x", io_vloadWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_245) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 11 and port 15 both writing to addr %x", io_vloadWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_246) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 11 and port 16 both writing to addr %x", io_vloadWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_247) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 11 and port 17 both writing to addr %x", io_vloadWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_248) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 11 and port 18 both writing to addr %x", io_vloadWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_249) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 11 and port 19 both writing to addr %x", io_vloadWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_250) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 11 and port 20 both writing to addr %x", io_vloadWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_251) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 11 and port 21 both writing to addr %x", io_vloadWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_252) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 11 and port 22 both writing to addr %x", io_vloadWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_253) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 11 and port 23 both writing to addr %x", io_vloadWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_254) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 11 and port 24 both writing to addr %x", io_vloadWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_255) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 11 and port 25 both writing to addr %x", io_vloadWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_256) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 11 and port 26 both writing to addr %x", io_vloadWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_257) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 11 and port 27 both writing to addr %x", io_vloadWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_258) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 12 and port 13 both writing to addr %x", io_vloadWrites_1_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_259) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 12 and port 14 both writing to addr %x", io_vloadWrites_1_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_260) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 12 and port 15 both writing to addr %x", io_vloadWrites_1_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_261) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 12 and port 16 both writing to addr %x", io_vloadWrites_1_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_262) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 12 and port 17 both writing to addr %x", io_vloadWrites_1_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_263) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 12 and port 18 both writing to addr %x", io_vloadWrites_1_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_264) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 12 and port 19 both writing to addr %x", io_vloadWrites_1_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_265) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 12 and port 20 both writing to addr %x", io_vloadWrites_1_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_266) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 12 and port 21 both writing to addr %x", io_vloadWrites_1_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_267) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 12 and port 22 both writing to addr %x", io_vloadWrites_1_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_268) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 12 and port 23 both writing to addr %x", io_vloadWrites_1_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_269) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 12 and port 24 both writing to addr %x", io_vloadWrites_1_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_270) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 12 and port 25 both writing to addr %x", io_vloadWrites_1_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_271) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 12 and port 26 both writing to addr %x", io_vloadWrites_1_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_272) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 12 and port 27 both writing to addr %x", io_vloadWrites_1_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_273) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 13 and port 14 both writing to addr %x", io_vloadWrites_2_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_274) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 13 and port 15 both writing to addr %x", io_vloadWrites_2_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_275) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 13 and port 16 both writing to addr %x", io_vloadWrites_2_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_276) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 13 and port 17 both writing to addr %x", io_vloadWrites_2_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_277) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 13 and port 18 both writing to addr %x", io_vloadWrites_2_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_278) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 13 and port 19 both writing to addr %x", io_vloadWrites_2_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_279) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 13 and port 20 both writing to addr %x", io_vloadWrites_2_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_280) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 13 and port 21 both writing to addr %x", io_vloadWrites_2_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_281) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 13 and port 22 both writing to addr %x", io_vloadWrites_2_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_282) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 13 and port 23 both writing to addr %x", io_vloadWrites_2_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_283) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 13 and port 24 both writing to addr %x", io_vloadWrites_2_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_284) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 13 and port 25 both writing to addr %x", io_vloadWrites_2_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_285) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 13 and port 26 both writing to addr %x", io_vloadWrites_2_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_286) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 13 and port 27 both writing to addr %x", io_vloadWrites_2_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_287) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 14 and port 15 both writing to addr %x", io_vloadWrites_3_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_288) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 14 and port 16 both writing to addr %x", io_vloadWrites_3_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_289) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 14 and port 17 both writing to addr %x", io_vloadWrites_3_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_290) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 14 and port 18 both writing to addr %x", io_vloadWrites_3_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_291) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 14 and port 19 both writing to addr %x", io_vloadWrites_3_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_292) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 14 and port 20 both writing to addr %x", io_vloadWrites_3_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_293) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 14 and port 21 both writing to addr %x", io_vloadWrites_3_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_294) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 14 and port 22 both writing to addr %x", io_vloadWrites_3_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_295) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 14 and port 23 both writing to addr %x", io_vloadWrites_3_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_296) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 14 and port 24 both writing to addr %x", io_vloadWrites_3_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_297) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 14 and port 25 both writing to addr %x", io_vloadWrites_3_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_298) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 14 and port 26 both writing to addr %x", io_vloadWrites_3_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_299) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 14 and port 27 both writing to addr %x", io_vloadWrites_3_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_300) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 15 and port 16 both writing to addr %x", io_vloadWrites_4_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_301) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 15 and port 17 both writing to addr %x", io_vloadWrites_4_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_302) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 15 and port 18 both writing to addr %x", io_vloadWrites_4_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_303) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 15 and port 19 both writing to addr %x", io_vloadWrites_4_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_304) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 15 and port 20 both writing to addr %x", io_vloadWrites_4_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_305) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 15 and port 21 both writing to addr %x", io_vloadWrites_4_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_306) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 15 and port 22 both writing to addr %x", io_vloadWrites_4_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_307) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 15 and port 23 both writing to addr %x", io_vloadWrites_4_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_308) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 15 and port 24 both writing to addr %x", io_vloadWrites_4_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_309) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 15 and port 25 both writing to addr %x", io_vloadWrites_4_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_310) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 15 and port 26 both writing to addr %x", io_vloadWrites_4_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_311) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 15 and port 27 both writing to addr %x", io_vloadWrites_4_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_312) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 16 and port 17 both writing to addr %x", io_vloadWrites_5_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_313) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 16 and port 18 both writing to addr %x", io_vloadWrites_5_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_314) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 16 and port 19 both writing to addr %x", io_vloadWrites_5_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_315) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 16 and port 20 both writing to addr %x", io_vloadWrites_5_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_316) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 16 and port 21 both writing to addr %x", io_vloadWrites_5_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_317) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 16 and port 22 both writing to addr %x", io_vloadWrites_5_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_318) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 16 and port 23 both writing to addr %x", io_vloadWrites_5_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_319) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 16 and port 24 both writing to addr %x", io_vloadWrites_5_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_320) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 16 and port 25 both writing to addr %x", io_vloadWrites_5_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_321) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 16 and port 26 both writing to addr %x", io_vloadWrites_5_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_322) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 16 and port 27 both writing to addr %x", io_vloadWrites_5_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_323) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 17 and port 18 both writing to addr %x", io_vloadWrites_6_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_324) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 17 and port 19 both writing to addr %x", io_vloadWrites_6_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_325) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 17 and port 20 both writing to addr %x", io_vloadWrites_6_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_326) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 17 and port 21 both writing to addr %x", io_vloadWrites_6_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_327) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 17 and port 22 both writing to addr %x", io_vloadWrites_6_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_328) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 17 and port 23 both writing to addr %x", io_vloadWrites_6_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_329) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 17 and port 24 both writing to addr %x", io_vloadWrites_6_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_330) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 17 and port 25 both writing to addr %x", io_vloadWrites_6_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_331) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 17 and port 26 both writing to addr %x", io_vloadWrites_6_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_332) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 17 and port 27 both writing to addr %x", io_vloadWrites_6_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_333) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 18 and port 19 both writing to addr %x", io_vloadWrites_7_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_334) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 18 and port 20 both writing to addr %x", io_vloadWrites_7_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_335) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 18 and port 21 both writing to addr %x", io_vloadWrites_7_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_336) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 18 and port 22 both writing to addr %x", io_vloadWrites_7_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_337) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 18 and port 23 both writing to addr %x", io_vloadWrites_7_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_338) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 18 and port 24 both writing to addr %x", io_vloadWrites_7_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_339) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 18 and port 25 both writing to addr %x", io_vloadWrites_7_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_340) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 18 and port 26 both writing to addr %x", io_vloadWrites_7_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_341) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 18 and port 27 both writing to addr %x", io_vloadWrites_7_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_342) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 19 and port 20 both writing to addr %x", io_flowScalarWrite_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_343) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 19 and port 21 both writing to addr %x", io_flowScalarWrite_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_344) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 19 and port 22 both writing to addr %x", io_flowScalarWrite_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_345) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 19 and port 23 both writing to addr %x", io_flowScalarWrite_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_346) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 19 and port 24 both writing to addr %x", io_flowScalarWrite_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_347) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 19 and port 25 both writing to addr %x", io_flowScalarWrite_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_348) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 19 and port 26 both writing to addr %x", io_flowScalarWrite_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_349) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 19 and port 27 both writing to addr %x", io_flowScalarWrite_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_350) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 20 and port 21 both writing to addr %x", io_flowVectorWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_351) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 20 and port 22 both writing to addr %x", io_flowVectorWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_352) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 20 and port 23 both writing to addr %x", io_flowVectorWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_353) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 20 and port 24 both writing to addr %x", io_flowVectorWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_354) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 20 and port 25 both writing to addr %x", io_flowVectorWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_355) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 20 and port 26 both writing to addr %x", io_flowVectorWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_356) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 20 and port 27 both writing to addr %x", io_flowVectorWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_357) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 21 and port 22 both writing to addr %x", io_flowVectorWrites_1_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_358) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 21 and port 23 both writing to addr %x", io_flowVectorWrites_1_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_359) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 21 and port 24 both writing to addr %x", io_flowVectorWrites_1_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_360) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 21 and port 25 both writing to addr %x", io_flowVectorWrites_1_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_361) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 21 and port 26 both writing to addr %x", io_flowVectorWrites_1_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_362) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 21 and port 27 both writing to addr %x", io_flowVectorWrites_1_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_363) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 22 and port 23 both writing to addr %x", io_flowVectorWrites_2_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_364) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 22 and port 24 both writing to addr %x", io_flowVectorWrites_2_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_365) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 22 and port 25 both writing to addr %x", io_flowVectorWrites_2_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_366) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 22 and port 26 both writing to addr %x", io_flowVectorWrites_2_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_367) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 22 and port 27 both writing to addr %x", io_flowVectorWrites_2_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_368) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 23 and port 24 both writing to addr %x", io_flowVectorWrites_3_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_369) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 23 and port 25 both writing to addr %x", io_flowVectorWrites_3_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_370) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 23 and port 26 both writing to addr %x", io_flowVectorWrites_3_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_371) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 23 and port 27 both writing to addr %x", io_flowVectorWrites_3_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_372) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 24 and port 25 both writing to addr %x", io_flowVectorWrites_4_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_373) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 24 and port 26 both writing to addr %x", io_flowVectorWrites_4_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_374) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 24 and port 27 both writing to addr %x", io_flowVectorWrites_4_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_375) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 25 and port 26 both writing to addr %x", io_flowVectorWrites_5_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_376) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 25 and port 27 both writing to addr %x", io_flowVectorWrites_5_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l84_377) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 26 and port 27 both writing to addr %x", io_flowVectorWrites_6_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
    end
  end


endmodule

module MemoryEngine (
  input  wire          io_loadSlots_0_valid,
  input  wire [2:0]    io_loadSlots_0_opcode,
  input  wire [10:0]   io_loadSlots_0_dest,
  input  wire [10:0]   io_loadSlots_0_addrReg,
  input  wire [2:0]    io_loadSlots_0_offset,
  input  wire [31:0]   io_loadSlots_0_immediate,
  input  wire          io_storeSlots_0_valid,
  input  wire [1:0]    io_storeSlots_0_opcode,
  input  wire [10:0]   io_storeSlots_0_addrReg,
  input  wire [10:0]   io_storeSlots_0_srcReg,
  input  wire          io_valid,
  input  wire [31:0]   io_loadAddrData_0,
  input  wire [31:0]   io_storeAddrData_0,
  input  wire [31:0]   io_storeSrcData_0,
  input  wire [31:0]   io_vstoreSrcData_0_0,
  input  wire [31:0]   io_vstoreSrcData_0_1,
  input  wire [31:0]   io_vstoreSrcData_0_2,
  input  wire [31:0]   io_vstoreSrcData_0_3,
  input  wire [31:0]   io_vstoreSrcData_0_4,
  input  wire [31:0]   io_vstoreSrcData_0_5,
  input  wire [31:0]   io_vstoreSrcData_0_6,
  input  wire [31:0]   io_vstoreSrcData_0_7,
  output reg           io_axiMaster_aw_valid,
  input  wire          io_axiMaster_aw_ready,
  output reg  [31:0]   io_axiMaster_aw_payload_addr,
  output wire [3:0]    io_axiMaster_aw_payload_id,
  output reg  [7:0]    io_axiMaster_aw_payload_len,
  output wire [2:0]    io_axiMaster_aw_payload_size,
  output wire [1:0]    io_axiMaster_aw_payload_burst,
  output reg           io_axiMaster_w_valid,
  input  wire          io_axiMaster_w_ready,
  output reg  [31:0]   io_axiMaster_w_payload_data,
  output wire [3:0]    io_axiMaster_w_payload_strb,
  output reg           io_axiMaster_w_payload_last,
  input  wire          io_axiMaster_b_valid,
  output wire          io_axiMaster_b_ready,
  input  wire [3:0]    io_axiMaster_b_payload_id,
  input  wire [1:0]    io_axiMaster_b_payload_resp,
  output reg           io_axiMaster_ar_valid,
  input  wire          io_axiMaster_ar_ready,
  output reg  [31:0]   io_axiMaster_ar_payload_addr,
  output wire [3:0]    io_axiMaster_ar_payload_id,
  output reg  [7:0]    io_axiMaster_ar_payload_len,
  output wire [2:0]    io_axiMaster_ar_payload_size,
  output wire [1:0]    io_axiMaster_ar_payload_burst,
  input  wire          io_axiMaster_r_valid,
  output wire          io_axiMaster_r_ready,
  input  wire [31:0]   io_axiMaster_r_payload_data,
  input  wire [3:0]    io_axiMaster_r_payload_id,
  input  wire [1:0]    io_axiMaster_r_payload_resp,
  input  wire          io_axiMaster_r_payload_last,
  output reg           io_loadWriteReqs_0_valid,
  output reg  [10:0]   io_loadWriteReqs_0_payload_addr,
  output reg  [31:0]   io_loadWriteReqs_0_payload_data,
  output reg           io_constWriteReqs_0_valid,
  output reg  [10:0]   io_constWriteReqs_0_payload_addr,
  output reg  [31:0]   io_constWriteReqs_0_payload_data,
  output reg           io_vloadWriteReqs_0_0_valid,
  output reg  [10:0]   io_vloadWriteReqs_0_0_payload_addr,
  output reg  [31:0]   io_vloadWriteReqs_0_0_payload_data,
  output reg           io_vloadWriteReqs_0_1_valid,
  output reg  [10:0]   io_vloadWriteReqs_0_1_payload_addr,
  output reg  [31:0]   io_vloadWriteReqs_0_1_payload_data,
  output reg           io_vloadWriteReqs_0_2_valid,
  output reg  [10:0]   io_vloadWriteReqs_0_2_payload_addr,
  output reg  [31:0]   io_vloadWriteReqs_0_2_payload_data,
  output reg           io_vloadWriteReqs_0_3_valid,
  output reg  [10:0]   io_vloadWriteReqs_0_3_payload_addr,
  output reg  [31:0]   io_vloadWriteReqs_0_3_payload_data,
  output reg           io_vloadWriteReqs_0_4_valid,
  output reg  [10:0]   io_vloadWriteReqs_0_4_payload_addr,
  output reg  [31:0]   io_vloadWriteReqs_0_4_payload_data,
  output reg           io_vloadWriteReqs_0_5_valid,
  output reg  [10:0]   io_vloadWriteReqs_0_5_payload_addr,
  output reg  [31:0]   io_vloadWriteReqs_0_5_payload_data,
  output reg           io_vloadWriteReqs_0_6_valid,
  output reg  [10:0]   io_vloadWriteReqs_0_6_payload_addr,
  output reg  [31:0]   io_vloadWriteReqs_0_6_payload_data,
  output reg           io_vloadWriteReqs_0_7_valid,
  output reg  [10:0]   io_vloadWriteReqs_0_7_payload_addr,
  output reg  [31:0]   io_vloadWriteReqs_0_7_payload_data,
  output reg           io_stall,
  input  wire          clk,
  input  wire          reset
);
  localparam MemState_IDLE = 4'd0;
  localparam MemState_LOAD_AR = 4'd1;
  localparam MemState_LOAD_R = 4'd2;
  localparam MemState_VLOAD_AR = 4'd3;
  localparam MemState_VLOAD_R = 4'd4;
  localparam MemState_STORE_AW = 4'd5;
  localparam MemState_STORE_W = 4'd6;
  localparam MemState_STORE_B = 4'd7;
  localparam MemState_VSTORE_AW = 4'd8;
  localparam MemState_VSTORE_W = 4'd9;
  localparam MemState_VSTORE_B = 4'd10;

  wire       [33:0]   _zz_capAddr;
  wire       [10:0]   _zz_capDest;
  wire       [33:0]   _zz_capAddr_1;
  wire       [31:0]   _zz_capAddr_2;
  wire       [31:0]   _zz_capAddr_3;
  wire       [33:0]   _zz_capAddr_4;
  wire       [33:0]   _zz_capAddr_5;
  wire       [33:0]   _zz_capAddr_6;
  reg        [3:0]    state;
  wire       [0:0]    slotIdx;
  reg        [3:0]    beatCount;
  wire                isStore;
  reg        [10:0]   capDest;
  reg        [31:0]   capAddr;
  reg        [2:0]    capOffset;
  reg        [0:0]    capSlotIdx;
  reg                 anyMemOp;
  wire                pendingLoads_0;
  wire                pendingStores_0;
  wire                when_MemoryEngine_l146;
  wire                when_MemoryEngine_l155;
  wire                when_MemoryEngine_l161;
  wire                when_MemoryEngine_l169;
  wire                when_MemoryEngine_l182;
  wire                when_MemoryEngine_l219;
  wire                when_MemoryEngine_l265;
  wire                when_MemoryEngine_l288;
  wire                when_MemoryEngine_l290;
  wire                when_MemoryEngine_l290_1;
  wire                when_MemoryEngine_l290_2;
  wire                when_MemoryEngine_l290_3;
  wire                when_MemoryEngine_l290_4;
  wire                when_MemoryEngine_l290_5;
  wire                when_MemoryEngine_l290_6;
  wire                when_MemoryEngine_l290_7;
  wire                when_MemoryEngine_l319;
  wire                when_MemoryEngine_l349;
  wire                when_MemoryEngine_l351;
  wire                when_MemoryEngine_l351_1;
  wire                when_MemoryEngine_l351_2;
  wire                when_MemoryEngine_l351_3;
  wire                when_MemoryEngine_l351_4;
  wire                when_MemoryEngine_l351_5;
  wire                when_MemoryEngine_l351_6;
  wire                when_MemoryEngine_l351_7;
  wire                when_MemoryEngine_l359;
  `ifndef SYNTHESIS
  reg [71:0] state_string;
  `endif


  assign _zz_capAddr = ({2'd0,io_loadAddrData_0} <<< 2'd2);
  assign _zz_capDest = {8'd0, io_loadSlots_0_offset};
  assign _zz_capAddr_1 = ({2'd0,_zz_capAddr_2} <<< 2'd2);
  assign _zz_capAddr_2 = (io_loadAddrData_0 + _zz_capAddr_3);
  assign _zz_capAddr_3 = {29'd0, io_loadSlots_0_offset};
  assign _zz_capAddr_4 = ({2'd0,io_loadAddrData_0} <<< 2'd2);
  assign _zz_capAddr_5 = ({2'd0,io_storeAddrData_0} <<< 2'd2);
  assign _zz_capAddr_6 = ({2'd0,io_storeAddrData_0} <<< 2'd2);
  `ifndef SYNTHESIS
  always @(*) begin
    case(state)
      MemState_IDLE : state_string = "IDLE     ";
      MemState_LOAD_AR : state_string = "LOAD_AR  ";
      MemState_LOAD_R : state_string = "LOAD_R   ";
      MemState_VLOAD_AR : state_string = "VLOAD_AR ";
      MemState_VLOAD_R : state_string = "VLOAD_R  ";
      MemState_STORE_AW : state_string = "STORE_AW ";
      MemState_STORE_W : state_string = "STORE_W  ";
      MemState_STORE_B : state_string = "STORE_B  ";
      MemState_VSTORE_AW : state_string = "VSTORE_AW";
      MemState_VSTORE_W : state_string = "VSTORE_W ";
      MemState_VSTORE_B : state_string = "VSTORE_B ";
      default : state_string = "?????????";
    endcase
  end
  `endif

  always @(*) begin
    io_stall = 1'b0;
    if(when_MemoryEngine_l169) begin
      io_stall = ((state != MemState_IDLE) || anyMemOp);
    end
  end

  always @(*) begin
    io_loadWriteReqs_0_valid = 1'b0;
    case(state)
      MemState_IDLE : begin
      end
      MemState_LOAD_AR : begin
      end
      MemState_LOAD_R : begin
        if(io_axiMaster_r_valid) begin
          if(when_MemoryEngine_l265) begin
            io_loadWriteReqs_0_valid = 1'b1;
          end
        end
      end
      MemState_VLOAD_AR : begin
      end
      MemState_VLOAD_R : begin
      end
      MemState_STORE_AW : begin
      end
      MemState_STORE_W : begin
      end
      MemState_STORE_B : begin
      end
      MemState_VSTORE_AW : begin
      end
      MemState_VSTORE_W : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_loadWriteReqs_0_payload_addr = 11'h0;
    case(state)
      MemState_IDLE : begin
      end
      MemState_LOAD_AR : begin
      end
      MemState_LOAD_R : begin
        if(io_axiMaster_r_valid) begin
          if(when_MemoryEngine_l265) begin
            io_loadWriteReqs_0_payload_addr = capDest;
          end
        end
      end
      MemState_VLOAD_AR : begin
      end
      MemState_VLOAD_R : begin
      end
      MemState_STORE_AW : begin
      end
      MemState_STORE_W : begin
      end
      MemState_STORE_B : begin
      end
      MemState_VSTORE_AW : begin
      end
      MemState_VSTORE_W : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_loadWriteReqs_0_payload_data = 32'h0;
    case(state)
      MemState_IDLE : begin
      end
      MemState_LOAD_AR : begin
      end
      MemState_LOAD_R : begin
        if(io_axiMaster_r_valid) begin
          if(when_MemoryEngine_l265) begin
            io_loadWriteReqs_0_payload_data = io_axiMaster_r_payload_data;
          end
        end
      end
      MemState_VLOAD_AR : begin
      end
      MemState_VLOAD_R : begin
      end
      MemState_STORE_AW : begin
      end
      MemState_STORE_W : begin
      end
      MemState_STORE_B : begin
      end
      MemState_VSTORE_AW : begin
      end
      MemState_VSTORE_W : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_constWriteReqs_0_valid = 1'b0;
    if(when_MemoryEngine_l161) begin
      io_constWriteReqs_0_valid = 1'b1;
    end
  end

  always @(*) begin
    io_constWriteReqs_0_payload_addr = 11'h0;
    if(when_MemoryEngine_l161) begin
      io_constWriteReqs_0_payload_addr = io_loadSlots_0_dest;
    end
  end

  always @(*) begin
    io_constWriteReqs_0_payload_data = 32'h0;
    if(when_MemoryEngine_l161) begin
      io_constWriteReqs_0_payload_data = io_loadSlots_0_immediate;
    end
  end

  always @(*) begin
    io_vloadWriteReqs_0_0_valid = 1'b0;
    case(state)
      MemState_IDLE : begin
      end
      MemState_LOAD_AR : begin
      end
      MemState_LOAD_R : begin
      end
      MemState_VLOAD_AR : begin
      end
      MemState_VLOAD_R : begin
        if(io_axiMaster_r_valid) begin
          if(when_MemoryEngine_l288) begin
            if(when_MemoryEngine_l290) begin
              io_vloadWriteReqs_0_0_valid = 1'b1;
            end
          end
        end
      end
      MemState_STORE_AW : begin
      end
      MemState_STORE_W : begin
      end
      MemState_STORE_B : begin
      end
      MemState_VSTORE_AW : begin
      end
      MemState_VSTORE_W : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_vloadWriteReqs_0_0_payload_addr = 11'h0;
    case(state)
      MemState_IDLE : begin
      end
      MemState_LOAD_AR : begin
      end
      MemState_LOAD_R : begin
      end
      MemState_VLOAD_AR : begin
      end
      MemState_VLOAD_R : begin
        if(io_axiMaster_r_valid) begin
          if(when_MemoryEngine_l288) begin
            if(when_MemoryEngine_l290) begin
              io_vloadWriteReqs_0_0_payload_addr = (capDest + 11'h0);
            end
          end
        end
      end
      MemState_STORE_AW : begin
      end
      MemState_STORE_W : begin
      end
      MemState_STORE_B : begin
      end
      MemState_VSTORE_AW : begin
      end
      MemState_VSTORE_W : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_vloadWriteReqs_0_0_payload_data = 32'h0;
    case(state)
      MemState_IDLE : begin
      end
      MemState_LOAD_AR : begin
      end
      MemState_LOAD_R : begin
      end
      MemState_VLOAD_AR : begin
      end
      MemState_VLOAD_R : begin
        if(io_axiMaster_r_valid) begin
          if(when_MemoryEngine_l288) begin
            if(when_MemoryEngine_l290) begin
              io_vloadWriteReqs_0_0_payload_data = io_axiMaster_r_payload_data;
            end
          end
        end
      end
      MemState_STORE_AW : begin
      end
      MemState_STORE_W : begin
      end
      MemState_STORE_B : begin
      end
      MemState_VSTORE_AW : begin
      end
      MemState_VSTORE_W : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_vloadWriteReqs_0_1_valid = 1'b0;
    case(state)
      MemState_IDLE : begin
      end
      MemState_LOAD_AR : begin
      end
      MemState_LOAD_R : begin
      end
      MemState_VLOAD_AR : begin
      end
      MemState_VLOAD_R : begin
        if(io_axiMaster_r_valid) begin
          if(when_MemoryEngine_l288) begin
            if(when_MemoryEngine_l290_1) begin
              io_vloadWriteReqs_0_1_valid = 1'b1;
            end
          end
        end
      end
      MemState_STORE_AW : begin
      end
      MemState_STORE_W : begin
      end
      MemState_STORE_B : begin
      end
      MemState_VSTORE_AW : begin
      end
      MemState_VSTORE_W : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_vloadWriteReqs_0_1_payload_addr = 11'h0;
    case(state)
      MemState_IDLE : begin
      end
      MemState_LOAD_AR : begin
      end
      MemState_LOAD_R : begin
      end
      MemState_VLOAD_AR : begin
      end
      MemState_VLOAD_R : begin
        if(io_axiMaster_r_valid) begin
          if(when_MemoryEngine_l288) begin
            if(when_MemoryEngine_l290_1) begin
              io_vloadWriteReqs_0_1_payload_addr = (capDest + 11'h001);
            end
          end
        end
      end
      MemState_STORE_AW : begin
      end
      MemState_STORE_W : begin
      end
      MemState_STORE_B : begin
      end
      MemState_VSTORE_AW : begin
      end
      MemState_VSTORE_W : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_vloadWriteReqs_0_1_payload_data = 32'h0;
    case(state)
      MemState_IDLE : begin
      end
      MemState_LOAD_AR : begin
      end
      MemState_LOAD_R : begin
      end
      MemState_VLOAD_AR : begin
      end
      MemState_VLOAD_R : begin
        if(io_axiMaster_r_valid) begin
          if(when_MemoryEngine_l288) begin
            if(when_MemoryEngine_l290_1) begin
              io_vloadWriteReqs_0_1_payload_data = io_axiMaster_r_payload_data;
            end
          end
        end
      end
      MemState_STORE_AW : begin
      end
      MemState_STORE_W : begin
      end
      MemState_STORE_B : begin
      end
      MemState_VSTORE_AW : begin
      end
      MemState_VSTORE_W : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_vloadWriteReqs_0_2_valid = 1'b0;
    case(state)
      MemState_IDLE : begin
      end
      MemState_LOAD_AR : begin
      end
      MemState_LOAD_R : begin
      end
      MemState_VLOAD_AR : begin
      end
      MemState_VLOAD_R : begin
        if(io_axiMaster_r_valid) begin
          if(when_MemoryEngine_l288) begin
            if(when_MemoryEngine_l290_2) begin
              io_vloadWriteReqs_0_2_valid = 1'b1;
            end
          end
        end
      end
      MemState_STORE_AW : begin
      end
      MemState_STORE_W : begin
      end
      MemState_STORE_B : begin
      end
      MemState_VSTORE_AW : begin
      end
      MemState_VSTORE_W : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_vloadWriteReqs_0_2_payload_addr = 11'h0;
    case(state)
      MemState_IDLE : begin
      end
      MemState_LOAD_AR : begin
      end
      MemState_LOAD_R : begin
      end
      MemState_VLOAD_AR : begin
      end
      MemState_VLOAD_R : begin
        if(io_axiMaster_r_valid) begin
          if(when_MemoryEngine_l288) begin
            if(when_MemoryEngine_l290_2) begin
              io_vloadWriteReqs_0_2_payload_addr = (capDest + 11'h002);
            end
          end
        end
      end
      MemState_STORE_AW : begin
      end
      MemState_STORE_W : begin
      end
      MemState_STORE_B : begin
      end
      MemState_VSTORE_AW : begin
      end
      MemState_VSTORE_W : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_vloadWriteReqs_0_2_payload_data = 32'h0;
    case(state)
      MemState_IDLE : begin
      end
      MemState_LOAD_AR : begin
      end
      MemState_LOAD_R : begin
      end
      MemState_VLOAD_AR : begin
      end
      MemState_VLOAD_R : begin
        if(io_axiMaster_r_valid) begin
          if(when_MemoryEngine_l288) begin
            if(when_MemoryEngine_l290_2) begin
              io_vloadWriteReqs_0_2_payload_data = io_axiMaster_r_payload_data;
            end
          end
        end
      end
      MemState_STORE_AW : begin
      end
      MemState_STORE_W : begin
      end
      MemState_STORE_B : begin
      end
      MemState_VSTORE_AW : begin
      end
      MemState_VSTORE_W : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_vloadWriteReqs_0_3_valid = 1'b0;
    case(state)
      MemState_IDLE : begin
      end
      MemState_LOAD_AR : begin
      end
      MemState_LOAD_R : begin
      end
      MemState_VLOAD_AR : begin
      end
      MemState_VLOAD_R : begin
        if(io_axiMaster_r_valid) begin
          if(when_MemoryEngine_l288) begin
            if(when_MemoryEngine_l290_3) begin
              io_vloadWriteReqs_0_3_valid = 1'b1;
            end
          end
        end
      end
      MemState_STORE_AW : begin
      end
      MemState_STORE_W : begin
      end
      MemState_STORE_B : begin
      end
      MemState_VSTORE_AW : begin
      end
      MemState_VSTORE_W : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_vloadWriteReqs_0_3_payload_addr = 11'h0;
    case(state)
      MemState_IDLE : begin
      end
      MemState_LOAD_AR : begin
      end
      MemState_LOAD_R : begin
      end
      MemState_VLOAD_AR : begin
      end
      MemState_VLOAD_R : begin
        if(io_axiMaster_r_valid) begin
          if(when_MemoryEngine_l288) begin
            if(when_MemoryEngine_l290_3) begin
              io_vloadWriteReqs_0_3_payload_addr = (capDest + 11'h003);
            end
          end
        end
      end
      MemState_STORE_AW : begin
      end
      MemState_STORE_W : begin
      end
      MemState_STORE_B : begin
      end
      MemState_VSTORE_AW : begin
      end
      MemState_VSTORE_W : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_vloadWriteReqs_0_3_payload_data = 32'h0;
    case(state)
      MemState_IDLE : begin
      end
      MemState_LOAD_AR : begin
      end
      MemState_LOAD_R : begin
      end
      MemState_VLOAD_AR : begin
      end
      MemState_VLOAD_R : begin
        if(io_axiMaster_r_valid) begin
          if(when_MemoryEngine_l288) begin
            if(when_MemoryEngine_l290_3) begin
              io_vloadWriteReqs_0_3_payload_data = io_axiMaster_r_payload_data;
            end
          end
        end
      end
      MemState_STORE_AW : begin
      end
      MemState_STORE_W : begin
      end
      MemState_STORE_B : begin
      end
      MemState_VSTORE_AW : begin
      end
      MemState_VSTORE_W : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_vloadWriteReqs_0_4_valid = 1'b0;
    case(state)
      MemState_IDLE : begin
      end
      MemState_LOAD_AR : begin
      end
      MemState_LOAD_R : begin
      end
      MemState_VLOAD_AR : begin
      end
      MemState_VLOAD_R : begin
        if(io_axiMaster_r_valid) begin
          if(when_MemoryEngine_l288) begin
            if(when_MemoryEngine_l290_4) begin
              io_vloadWriteReqs_0_4_valid = 1'b1;
            end
          end
        end
      end
      MemState_STORE_AW : begin
      end
      MemState_STORE_W : begin
      end
      MemState_STORE_B : begin
      end
      MemState_VSTORE_AW : begin
      end
      MemState_VSTORE_W : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_vloadWriteReqs_0_4_payload_addr = 11'h0;
    case(state)
      MemState_IDLE : begin
      end
      MemState_LOAD_AR : begin
      end
      MemState_LOAD_R : begin
      end
      MemState_VLOAD_AR : begin
      end
      MemState_VLOAD_R : begin
        if(io_axiMaster_r_valid) begin
          if(when_MemoryEngine_l288) begin
            if(when_MemoryEngine_l290_4) begin
              io_vloadWriteReqs_0_4_payload_addr = (capDest + 11'h004);
            end
          end
        end
      end
      MemState_STORE_AW : begin
      end
      MemState_STORE_W : begin
      end
      MemState_STORE_B : begin
      end
      MemState_VSTORE_AW : begin
      end
      MemState_VSTORE_W : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_vloadWriteReqs_0_4_payload_data = 32'h0;
    case(state)
      MemState_IDLE : begin
      end
      MemState_LOAD_AR : begin
      end
      MemState_LOAD_R : begin
      end
      MemState_VLOAD_AR : begin
      end
      MemState_VLOAD_R : begin
        if(io_axiMaster_r_valid) begin
          if(when_MemoryEngine_l288) begin
            if(when_MemoryEngine_l290_4) begin
              io_vloadWriteReqs_0_4_payload_data = io_axiMaster_r_payload_data;
            end
          end
        end
      end
      MemState_STORE_AW : begin
      end
      MemState_STORE_W : begin
      end
      MemState_STORE_B : begin
      end
      MemState_VSTORE_AW : begin
      end
      MemState_VSTORE_W : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_vloadWriteReqs_0_5_valid = 1'b0;
    case(state)
      MemState_IDLE : begin
      end
      MemState_LOAD_AR : begin
      end
      MemState_LOAD_R : begin
      end
      MemState_VLOAD_AR : begin
      end
      MemState_VLOAD_R : begin
        if(io_axiMaster_r_valid) begin
          if(when_MemoryEngine_l288) begin
            if(when_MemoryEngine_l290_5) begin
              io_vloadWriteReqs_0_5_valid = 1'b1;
            end
          end
        end
      end
      MemState_STORE_AW : begin
      end
      MemState_STORE_W : begin
      end
      MemState_STORE_B : begin
      end
      MemState_VSTORE_AW : begin
      end
      MemState_VSTORE_W : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_vloadWriteReqs_0_5_payload_addr = 11'h0;
    case(state)
      MemState_IDLE : begin
      end
      MemState_LOAD_AR : begin
      end
      MemState_LOAD_R : begin
      end
      MemState_VLOAD_AR : begin
      end
      MemState_VLOAD_R : begin
        if(io_axiMaster_r_valid) begin
          if(when_MemoryEngine_l288) begin
            if(when_MemoryEngine_l290_5) begin
              io_vloadWriteReqs_0_5_payload_addr = (capDest + 11'h005);
            end
          end
        end
      end
      MemState_STORE_AW : begin
      end
      MemState_STORE_W : begin
      end
      MemState_STORE_B : begin
      end
      MemState_VSTORE_AW : begin
      end
      MemState_VSTORE_W : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_vloadWriteReqs_0_5_payload_data = 32'h0;
    case(state)
      MemState_IDLE : begin
      end
      MemState_LOAD_AR : begin
      end
      MemState_LOAD_R : begin
      end
      MemState_VLOAD_AR : begin
      end
      MemState_VLOAD_R : begin
        if(io_axiMaster_r_valid) begin
          if(when_MemoryEngine_l288) begin
            if(when_MemoryEngine_l290_5) begin
              io_vloadWriteReqs_0_5_payload_data = io_axiMaster_r_payload_data;
            end
          end
        end
      end
      MemState_STORE_AW : begin
      end
      MemState_STORE_W : begin
      end
      MemState_STORE_B : begin
      end
      MemState_VSTORE_AW : begin
      end
      MemState_VSTORE_W : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_vloadWriteReqs_0_6_valid = 1'b0;
    case(state)
      MemState_IDLE : begin
      end
      MemState_LOAD_AR : begin
      end
      MemState_LOAD_R : begin
      end
      MemState_VLOAD_AR : begin
      end
      MemState_VLOAD_R : begin
        if(io_axiMaster_r_valid) begin
          if(when_MemoryEngine_l288) begin
            if(when_MemoryEngine_l290_6) begin
              io_vloadWriteReqs_0_6_valid = 1'b1;
            end
          end
        end
      end
      MemState_STORE_AW : begin
      end
      MemState_STORE_W : begin
      end
      MemState_STORE_B : begin
      end
      MemState_VSTORE_AW : begin
      end
      MemState_VSTORE_W : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_vloadWriteReqs_0_6_payload_addr = 11'h0;
    case(state)
      MemState_IDLE : begin
      end
      MemState_LOAD_AR : begin
      end
      MemState_LOAD_R : begin
      end
      MemState_VLOAD_AR : begin
      end
      MemState_VLOAD_R : begin
        if(io_axiMaster_r_valid) begin
          if(when_MemoryEngine_l288) begin
            if(when_MemoryEngine_l290_6) begin
              io_vloadWriteReqs_0_6_payload_addr = (capDest + 11'h006);
            end
          end
        end
      end
      MemState_STORE_AW : begin
      end
      MemState_STORE_W : begin
      end
      MemState_STORE_B : begin
      end
      MemState_VSTORE_AW : begin
      end
      MemState_VSTORE_W : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_vloadWriteReqs_0_6_payload_data = 32'h0;
    case(state)
      MemState_IDLE : begin
      end
      MemState_LOAD_AR : begin
      end
      MemState_LOAD_R : begin
      end
      MemState_VLOAD_AR : begin
      end
      MemState_VLOAD_R : begin
        if(io_axiMaster_r_valid) begin
          if(when_MemoryEngine_l288) begin
            if(when_MemoryEngine_l290_6) begin
              io_vloadWriteReqs_0_6_payload_data = io_axiMaster_r_payload_data;
            end
          end
        end
      end
      MemState_STORE_AW : begin
      end
      MemState_STORE_W : begin
      end
      MemState_STORE_B : begin
      end
      MemState_VSTORE_AW : begin
      end
      MemState_VSTORE_W : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_vloadWriteReqs_0_7_valid = 1'b0;
    case(state)
      MemState_IDLE : begin
      end
      MemState_LOAD_AR : begin
      end
      MemState_LOAD_R : begin
      end
      MemState_VLOAD_AR : begin
      end
      MemState_VLOAD_R : begin
        if(io_axiMaster_r_valid) begin
          if(when_MemoryEngine_l288) begin
            if(when_MemoryEngine_l290_7) begin
              io_vloadWriteReqs_0_7_valid = 1'b1;
            end
          end
        end
      end
      MemState_STORE_AW : begin
      end
      MemState_STORE_W : begin
      end
      MemState_STORE_B : begin
      end
      MemState_VSTORE_AW : begin
      end
      MemState_VSTORE_W : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_vloadWriteReqs_0_7_payload_addr = 11'h0;
    case(state)
      MemState_IDLE : begin
      end
      MemState_LOAD_AR : begin
      end
      MemState_LOAD_R : begin
      end
      MemState_VLOAD_AR : begin
      end
      MemState_VLOAD_R : begin
        if(io_axiMaster_r_valid) begin
          if(when_MemoryEngine_l288) begin
            if(when_MemoryEngine_l290_7) begin
              io_vloadWriteReqs_0_7_payload_addr = (capDest + 11'h007);
            end
          end
        end
      end
      MemState_STORE_AW : begin
      end
      MemState_STORE_W : begin
      end
      MemState_STORE_B : begin
      end
      MemState_VSTORE_AW : begin
      end
      MemState_VSTORE_W : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_vloadWriteReqs_0_7_payload_data = 32'h0;
    case(state)
      MemState_IDLE : begin
      end
      MemState_LOAD_AR : begin
      end
      MemState_LOAD_R : begin
      end
      MemState_VLOAD_AR : begin
      end
      MemState_VLOAD_R : begin
        if(io_axiMaster_r_valid) begin
          if(when_MemoryEngine_l288) begin
            if(when_MemoryEngine_l290_7) begin
              io_vloadWriteReqs_0_7_payload_data = io_axiMaster_r_payload_data;
            end
          end
        end
      end
      MemState_STORE_AW : begin
      end
      MemState_STORE_W : begin
      end
      MemState_STORE_B : begin
      end
      MemState_VSTORE_AW : begin
      end
      MemState_VSTORE_W : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_axiMaster_aw_valid = 1'b0;
    case(state)
      MemState_IDLE : begin
      end
      MemState_LOAD_AR : begin
      end
      MemState_LOAD_R : begin
      end
      MemState_VLOAD_AR : begin
      end
      MemState_VLOAD_R : begin
      end
      MemState_STORE_AW : begin
        io_axiMaster_aw_valid = 1'b1;
      end
      MemState_STORE_W : begin
      end
      MemState_STORE_B : begin
      end
      MemState_VSTORE_AW : begin
        io_axiMaster_aw_valid = 1'b1;
      end
      MemState_VSTORE_W : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_axiMaster_aw_payload_addr = 32'h0;
    case(state)
      MemState_IDLE : begin
      end
      MemState_LOAD_AR : begin
      end
      MemState_LOAD_R : begin
      end
      MemState_VLOAD_AR : begin
      end
      MemState_VLOAD_R : begin
      end
      MemState_STORE_AW : begin
        io_axiMaster_aw_payload_addr = capAddr;
      end
      MemState_STORE_W : begin
      end
      MemState_STORE_B : begin
      end
      MemState_VSTORE_AW : begin
        io_axiMaster_aw_payload_addr = capAddr;
      end
      MemState_VSTORE_W : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_axiMaster_aw_payload_len = 8'h0;
    case(state)
      MemState_IDLE : begin
      end
      MemState_LOAD_AR : begin
      end
      MemState_LOAD_R : begin
      end
      MemState_VLOAD_AR : begin
      end
      MemState_VLOAD_R : begin
      end
      MemState_STORE_AW : begin
        io_axiMaster_aw_payload_len = 8'h0;
      end
      MemState_STORE_W : begin
      end
      MemState_STORE_B : begin
      end
      MemState_VSTORE_AW : begin
        io_axiMaster_aw_payload_len = 8'h07;
      end
      MemState_VSTORE_W : begin
      end
      default : begin
      end
    endcase
  end

  assign io_axiMaster_aw_payload_size = 3'b010;
  assign io_axiMaster_aw_payload_burst = 2'b01;
  assign io_axiMaster_aw_payload_id = 4'b0000;
  always @(*) begin
    io_axiMaster_w_valid = 1'b0;
    case(state)
      MemState_IDLE : begin
      end
      MemState_LOAD_AR : begin
      end
      MemState_LOAD_R : begin
      end
      MemState_VLOAD_AR : begin
      end
      MemState_VLOAD_R : begin
      end
      MemState_STORE_AW : begin
      end
      MemState_STORE_W : begin
        io_axiMaster_w_valid = 1'b1;
      end
      MemState_STORE_B : begin
      end
      MemState_VSTORE_AW : begin
      end
      MemState_VSTORE_W : begin
        io_axiMaster_w_valid = 1'b1;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_axiMaster_w_payload_data = 32'h0;
    case(state)
      MemState_IDLE : begin
      end
      MemState_LOAD_AR : begin
      end
      MemState_LOAD_R : begin
      end
      MemState_VLOAD_AR : begin
      end
      MemState_VLOAD_R : begin
      end
      MemState_STORE_AW : begin
      end
      MemState_STORE_W : begin
        if(when_MemoryEngine_l319) begin
          io_axiMaster_w_payload_data = io_storeSrcData_0;
        end
      end
      MemState_STORE_B : begin
      end
      MemState_VSTORE_AW : begin
      end
      MemState_VSTORE_W : begin
        if(when_MemoryEngine_l349) begin
          if(when_MemoryEngine_l351) begin
            io_axiMaster_w_payload_data = io_vstoreSrcData_0_0;
          end
          if(when_MemoryEngine_l351_1) begin
            io_axiMaster_w_payload_data = io_vstoreSrcData_0_1;
          end
          if(when_MemoryEngine_l351_2) begin
            io_axiMaster_w_payload_data = io_vstoreSrcData_0_2;
          end
          if(when_MemoryEngine_l351_3) begin
            io_axiMaster_w_payload_data = io_vstoreSrcData_0_3;
          end
          if(when_MemoryEngine_l351_4) begin
            io_axiMaster_w_payload_data = io_vstoreSrcData_0_4;
          end
          if(when_MemoryEngine_l351_5) begin
            io_axiMaster_w_payload_data = io_vstoreSrcData_0_5;
          end
          if(when_MemoryEngine_l351_6) begin
            io_axiMaster_w_payload_data = io_vstoreSrcData_0_6;
          end
          if(when_MemoryEngine_l351_7) begin
            io_axiMaster_w_payload_data = io_vstoreSrcData_0_7;
          end
        end
      end
      default : begin
      end
    endcase
  end

  assign io_axiMaster_w_payload_strb = 4'b1111;
  always @(*) begin
    io_axiMaster_w_payload_last = 1'b1;
    case(state)
      MemState_IDLE : begin
      end
      MemState_LOAD_AR : begin
      end
      MemState_LOAD_R : begin
      end
      MemState_VLOAD_AR : begin
      end
      MemState_VLOAD_R : begin
      end
      MemState_STORE_AW : begin
      end
      MemState_STORE_W : begin
        io_axiMaster_w_payload_last = 1'b1;
      end
      MemState_STORE_B : begin
      end
      MemState_VSTORE_AW : begin
      end
      MemState_VSTORE_W : begin
        io_axiMaster_w_payload_last = (beatCount == 4'b0111);
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_axiMaster_ar_valid = 1'b0;
    case(state)
      MemState_IDLE : begin
      end
      MemState_LOAD_AR : begin
        io_axiMaster_ar_valid = 1'b1;
      end
      MemState_LOAD_R : begin
      end
      MemState_VLOAD_AR : begin
        io_axiMaster_ar_valid = 1'b1;
      end
      MemState_VLOAD_R : begin
      end
      MemState_STORE_AW : begin
      end
      MemState_STORE_W : begin
      end
      MemState_STORE_B : begin
      end
      MemState_VSTORE_AW : begin
      end
      MemState_VSTORE_W : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_axiMaster_ar_payload_addr = 32'h0;
    case(state)
      MemState_IDLE : begin
      end
      MemState_LOAD_AR : begin
        io_axiMaster_ar_payload_addr = capAddr;
      end
      MemState_LOAD_R : begin
      end
      MemState_VLOAD_AR : begin
        io_axiMaster_ar_payload_addr = capAddr;
      end
      MemState_VLOAD_R : begin
      end
      MemState_STORE_AW : begin
      end
      MemState_STORE_W : begin
      end
      MemState_STORE_B : begin
      end
      MemState_VSTORE_AW : begin
      end
      MemState_VSTORE_W : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_axiMaster_ar_payload_len = 8'h0;
    case(state)
      MemState_IDLE : begin
      end
      MemState_LOAD_AR : begin
        io_axiMaster_ar_payload_len = 8'h0;
      end
      MemState_LOAD_R : begin
      end
      MemState_VLOAD_AR : begin
        io_axiMaster_ar_payload_len = 8'h07;
      end
      MemState_VLOAD_R : begin
      end
      MemState_STORE_AW : begin
      end
      MemState_STORE_W : begin
      end
      MemState_STORE_B : begin
      end
      MemState_VSTORE_AW : begin
      end
      MemState_VSTORE_W : begin
      end
      default : begin
      end
    endcase
  end

  assign io_axiMaster_ar_payload_size = 3'b010;
  assign io_axiMaster_ar_payload_burst = 2'b01;
  assign io_axiMaster_ar_payload_id = 4'b0000;
  assign io_axiMaster_r_ready = 1'b1;
  assign io_axiMaster_b_ready = 1'b1;
  assign slotIdx = 1'b0;
  assign isStore = 1'b0;
  always @(*) begin
    anyMemOp = 1'b0;
    if(when_MemoryEngine_l146) begin
      anyMemOp = 1'b1;
    end
    if(when_MemoryEngine_l155) begin
      anyMemOp = 1'b1;
    end
  end

  assign when_MemoryEngine_l146 = ((io_loadSlots_0_valid && io_valid) && (((io_loadSlots_0_opcode == 3'b001) || (io_loadSlots_0_opcode == 3'b010)) || (io_loadSlots_0_opcode == 3'b011)));
  assign pendingLoads_0 = when_MemoryEngine_l146;
  assign when_MemoryEngine_l155 = ((io_storeSlots_0_valid && io_valid) && ((io_storeSlots_0_opcode == 2'b01) || (io_storeSlots_0_opcode == 2'b10)));
  assign pendingStores_0 = when_MemoryEngine_l155;
  assign when_MemoryEngine_l161 = ((io_loadSlots_0_valid && io_valid) && (io_loadSlots_0_opcode == 3'b100));
  assign when_MemoryEngine_l169 = ((state != MemState_IDLE) || anyMemOp);
  assign when_MemoryEngine_l182 = (|pendingLoads_0);
  assign when_MemoryEngine_l219 = (|pendingStores_0);
  assign when_MemoryEngine_l265 = (capSlotIdx == 1'b0);
  assign when_MemoryEngine_l288 = (capSlotIdx == 1'b0);
  assign when_MemoryEngine_l290 = (beatCount == 4'b0000);
  assign when_MemoryEngine_l290_1 = (beatCount == 4'b0001);
  assign when_MemoryEngine_l290_2 = (beatCount == 4'b0010);
  assign when_MemoryEngine_l290_3 = (beatCount == 4'b0011);
  assign when_MemoryEngine_l290_4 = (beatCount == 4'b0100);
  assign when_MemoryEngine_l290_5 = (beatCount == 4'b0101);
  assign when_MemoryEngine_l290_6 = (beatCount == 4'b0110);
  assign when_MemoryEngine_l290_7 = (beatCount == 4'b0111);
  assign when_MemoryEngine_l319 = (capSlotIdx == 1'b0);
  assign when_MemoryEngine_l349 = (capSlotIdx == 1'b0);
  assign when_MemoryEngine_l351 = (beatCount == 4'b0000);
  assign when_MemoryEngine_l351_1 = (beatCount == 4'b0001);
  assign when_MemoryEngine_l351_2 = (beatCount == 4'b0010);
  assign when_MemoryEngine_l351_3 = (beatCount == 4'b0011);
  assign when_MemoryEngine_l351_4 = (beatCount == 4'b0100);
  assign when_MemoryEngine_l351_5 = (beatCount == 4'b0101);
  assign when_MemoryEngine_l351_6 = (beatCount == 4'b0110);
  assign when_MemoryEngine_l351_7 = (beatCount == 4'b0111);
  assign when_MemoryEngine_l359 = (beatCount == 4'b0111);
  always @(posedge clk) begin
    if(reset) begin
      state <= MemState_IDLE;
      beatCount <= 4'b0000;
    end else begin
      case(state)
        MemState_IDLE : begin
          if(anyMemOp) begin
            if(when_MemoryEngine_l182) begin
              if(pendingLoads_0) begin
                case(io_loadSlots_0_opcode)
                  3'b001 : begin
                    state <= MemState_LOAD_AR;
                  end
                  3'b010 : begin
                    state <= MemState_LOAD_AR;
                  end
                  3'b011 : begin
                    beatCount <= 4'b0000;
                    state <= MemState_VLOAD_AR;
                  end
                  default : begin
                  end
                endcase
              end
            end else begin
              if(when_MemoryEngine_l219) begin
                if(pendingStores_0) begin
                  case(io_storeSlots_0_opcode)
                    2'b01 : begin
                      state <= MemState_STORE_AW;
                    end
                    2'b10 : begin
                      beatCount <= 4'b0000;
                      state <= MemState_VSTORE_AW;
                    end
                    default : begin
                    end
                  endcase
                end
              end
            end
          end
        end
        MemState_LOAD_AR : begin
          if(io_axiMaster_ar_ready) begin
            state <= MemState_LOAD_R;
          end
        end
        MemState_LOAD_R : begin
          if(io_axiMaster_r_valid) begin
            state <= MemState_IDLE;
          end
        end
        MemState_VLOAD_AR : begin
          if(io_axiMaster_ar_ready) begin
            state <= MemState_VLOAD_R;
          end
        end
        MemState_VLOAD_R : begin
          if(io_axiMaster_r_valid) begin
            beatCount <= (beatCount + 4'b0001);
            if(io_axiMaster_r_payload_last) begin
              state <= MemState_IDLE;
            end
          end
        end
        MemState_STORE_AW : begin
          if(io_axiMaster_aw_ready) begin
            state <= MemState_STORE_W;
          end
        end
        MemState_STORE_W : begin
          if(io_axiMaster_w_ready) begin
            state <= MemState_STORE_B;
          end
        end
        MemState_STORE_B : begin
          if(io_axiMaster_b_valid) begin
            state <= MemState_IDLE;
          end
        end
        MemState_VSTORE_AW : begin
          if(io_axiMaster_aw_ready) begin
            beatCount <= 4'b0000;
            state <= MemState_VSTORE_W;
          end
        end
        MemState_VSTORE_W : begin
          if(io_axiMaster_w_ready) begin
            beatCount <= (beatCount + 4'b0001);
            if(when_MemoryEngine_l359) begin
              state <= MemState_VSTORE_B;
            end
          end
        end
        default : begin
          if(io_axiMaster_b_valid) begin
            state <= MemState_IDLE;
          end
        end
      endcase
    end
  end

  always @(posedge clk) begin
    case(state)
      MemState_IDLE : begin
        if(anyMemOp) begin
          if(when_MemoryEngine_l182) begin
            if(pendingLoads_0) begin
              case(io_loadSlots_0_opcode)
                3'b001 : begin
                  capDest <= io_loadSlots_0_dest;
                  capAddr <= _zz_capAddr[31:0];
                  capSlotIdx <= 1'b0;
                end
                3'b010 : begin
                  capDest <= (io_loadSlots_0_dest + _zz_capDest);
                  capAddr <= _zz_capAddr_1[31:0];
                  capSlotIdx <= 1'b0;
                end
                3'b011 : begin
                  capDest <= io_loadSlots_0_dest;
                  capAddr <= _zz_capAddr_4[31:0];
                  capSlotIdx <= 1'b0;
                end
                default : begin
                end
              endcase
            end
          end else begin
            if(when_MemoryEngine_l219) begin
              if(pendingStores_0) begin
                case(io_storeSlots_0_opcode)
                  2'b01 : begin
                    capAddr <= _zz_capAddr_5[31:0];
                    capSlotIdx <= 1'b0;
                  end
                  2'b10 : begin
                    capAddr <= _zz_capAddr_6[31:0];
                    capSlotIdx <= 1'b0;
                  end
                  default : begin
                  end
                endcase
              end
            end
          end
        end
      end
      MemState_LOAD_AR : begin
      end
      MemState_LOAD_R : begin
      end
      MemState_VLOAD_AR : begin
      end
      MemState_VLOAD_R : begin
      end
      MemState_STORE_AW : begin
      end
      MemState_STORE_W : begin
      end
      MemState_STORE_B : begin
      end
      MemState_VSTORE_AW : begin
      end
      MemState_VSTORE_W : begin
      end
      default : begin
      end
    endcase
  end


endmodule

module FlowEngine (
  input  wire          io_slot_valid,
  input  wire [3:0]    io_slot_opcode,
  input  wire [10:0]   io_slot_dest,
  input  wire [10:0]   io_slot_operandA,
  input  wire [10:0]   io_slot_operandB,
  input  wire [9:0]    io_slot_immediate,
  input  wire          io_valid,
  input  wire [9:0]    io_currentPc,
  input  wire [31:0]   io_operandCond,
  input  wire [31:0]   io_operandA,
  input  wire [31:0]   io_operandB,
  input  wire [31:0]   io_vCond_0,
  input  wire [31:0]   io_vCond_1,
  input  wire [31:0]   io_vCond_2,
  input  wire [31:0]   io_vCond_3,
  input  wire [31:0]   io_vCond_4,
  input  wire [31:0]   io_vCond_5,
  input  wire [31:0]   io_vCond_6,
  input  wire [31:0]   io_vCond_7,
  input  wire [31:0]   io_vSrcA_0,
  input  wire [31:0]   io_vSrcA_1,
  input  wire [31:0]   io_vSrcA_2,
  input  wire [31:0]   io_vSrcA_3,
  input  wire [31:0]   io_vSrcA_4,
  input  wire [31:0]   io_vSrcA_5,
  input  wire [31:0]   io_vSrcA_6,
  input  wire [31:0]   io_vSrcA_7,
  input  wire [31:0]   io_vSrcB_0,
  input  wire [31:0]   io_vSrcB_1,
  input  wire [31:0]   io_vSrcB_2,
  input  wire [31:0]   io_vSrcB_3,
  input  wire [31:0]   io_vSrcB_4,
  input  wire [31:0]   io_vSrcB_5,
  input  wire [31:0]   io_vSrcB_6,
  input  wire [31:0]   io_vSrcB_7,
  output reg           io_scalarWriteReq_valid,
  output reg  [10:0]   io_scalarWriteReq_payload_addr,
  output reg  [31:0]   io_scalarWriteReq_payload_data,
  output reg           io_vectorWriteReqs_0_valid,
  output reg  [10:0]   io_vectorWriteReqs_0_payload_addr,
  output reg  [31:0]   io_vectorWriteReqs_0_payload_data,
  output reg           io_vectorWriteReqs_1_valid,
  output reg  [10:0]   io_vectorWriteReqs_1_payload_addr,
  output reg  [31:0]   io_vectorWriteReqs_1_payload_data,
  output reg           io_vectorWriteReqs_2_valid,
  output reg  [10:0]   io_vectorWriteReqs_2_payload_addr,
  output reg  [31:0]   io_vectorWriteReqs_2_payload_data,
  output reg           io_vectorWriteReqs_3_valid,
  output reg  [10:0]   io_vectorWriteReqs_3_payload_addr,
  output reg  [31:0]   io_vectorWriteReqs_3_payload_data,
  output reg           io_vectorWriteReqs_4_valid,
  output reg  [10:0]   io_vectorWriteReqs_4_payload_addr,
  output reg  [31:0]   io_vectorWriteReqs_4_payload_data,
  output reg           io_vectorWriteReqs_5_valid,
  output reg  [10:0]   io_vectorWriteReqs_5_payload_addr,
  output reg  [31:0]   io_vectorWriteReqs_5_payload_data,
  output reg           io_vectorWriteReqs_6_valid,
  output reg  [10:0]   io_vectorWriteReqs_6_payload_addr,
  output reg  [31:0]   io_vectorWriteReqs_6_payload_data,
  output reg           io_vectorWriteReqs_7_valid,
  output reg  [10:0]   io_vectorWriteReqs_7_payload_addr,
  output reg  [31:0]   io_vectorWriteReqs_7_payload_data,
  output reg           io_jumpTarget_valid,
  output reg  [9:0]    io_jumpTarget_payload,
  output reg           io_halt
);

  wire       [31:0]   _zz_io_scalarWriteReq_payload_data;
  wire       [9:0]    _zz_io_scalarWriteReq_payload_data_1;
  wire       [20:0]   _zz_io_jumpTarget_payload;
  wire       [9:0]    _zz_io_jumpTarget_payload_1;
  wire       [9:0]    _zz_io_jumpTarget_payload_2;
  wire       [9:0]    _zz_io_jumpTarget_payload_3;
  wire       [20:0]   _zz_io_jumpTarget_payload_4;
  wire                slotValid;
  wire                when_FlowEngine_l109;
  wire                when_FlowEngine_l118;

  assign _zz_io_scalarWriteReq_payload_data_1 = io_slot_immediate;
  assign _zz_io_scalarWriteReq_payload_data = {{22{_zz_io_scalarWriteReq_payload_data_1[9]}}, _zz_io_scalarWriteReq_payload_data_1};
  assign _zz_io_jumpTarget_payload = {io_slot_operandB,io_slot_immediate};
  assign _zz_io_jumpTarget_payload_1 = ($signed(_zz_io_jumpTarget_payload_2) + $signed(_zz_io_jumpTarget_payload_3));
  assign _zz_io_jumpTarget_payload_2 = io_currentPc;
  assign _zz_io_jumpTarget_payload_3 = io_slot_immediate;
  assign _zz_io_jumpTarget_payload_4 = {io_slot_operandB,io_slot_immediate};
  assign slotValid = (io_slot_valid && io_valid);
  always @(*) begin
    io_scalarWriteReq_valid = 1'b0;
    if(slotValid) begin
      case(io_slot_opcode)
        4'b0001 : begin
          io_scalarWriteReq_valid = 1'b1;
        end
        4'b0011 : begin
          io_scalarWriteReq_valid = 1'b1;
        end
        4'b1001 : begin
          io_scalarWriteReq_valid = 1'b1;
        end
        default : begin
        end
      endcase
    end
  end

  always @(*) begin
    io_scalarWriteReq_payload_addr = 11'h0;
    if(slotValid) begin
      case(io_slot_opcode)
        4'b0001 : begin
          io_scalarWriteReq_payload_addr = io_slot_dest;
        end
        4'b0011 : begin
          io_scalarWriteReq_payload_addr = io_slot_dest;
        end
        4'b1001 : begin
          io_scalarWriteReq_payload_addr = io_slot_dest;
        end
        default : begin
        end
      endcase
    end
  end

  always @(*) begin
    io_scalarWriteReq_payload_data = 32'h0;
    if(slotValid) begin
      case(io_slot_opcode)
        4'b0001 : begin
          io_scalarWriteReq_payload_data = ((io_operandCond != 32'h0) ? io_operandA : io_operandB);
        end
        4'b0011 : begin
          io_scalarWriteReq_payload_data = (io_operandCond + _zz_io_scalarWriteReq_payload_data);
        end
        4'b1001 : begin
          io_scalarWriteReq_payload_data = 32'h0;
        end
        default : begin
        end
      endcase
    end
  end

  always @(*) begin
    io_vectorWriteReqs_0_valid = 1'b0;
    if(slotValid) begin
      case(io_slot_opcode)
        4'b0010 : begin
          io_vectorWriteReqs_0_valid = 1'b1;
        end
        default : begin
        end
      endcase
    end
  end

  always @(*) begin
    io_vectorWriteReqs_0_payload_addr = 11'h0;
    if(slotValid) begin
      case(io_slot_opcode)
        4'b0010 : begin
          io_vectorWriteReqs_0_payload_addr = (io_slot_dest + 11'h0);
        end
        default : begin
        end
      endcase
    end
  end

  always @(*) begin
    io_vectorWriteReqs_0_payload_data = 32'h0;
    if(slotValid) begin
      case(io_slot_opcode)
        4'b0010 : begin
          io_vectorWriteReqs_0_payload_data = ((io_vCond_0 != 32'h0) ? io_vSrcA_0 : io_vSrcB_0);
        end
        default : begin
        end
      endcase
    end
  end

  always @(*) begin
    io_vectorWriteReqs_1_valid = 1'b0;
    if(slotValid) begin
      case(io_slot_opcode)
        4'b0010 : begin
          io_vectorWriteReqs_1_valid = 1'b1;
        end
        default : begin
        end
      endcase
    end
  end

  always @(*) begin
    io_vectorWriteReqs_1_payload_addr = 11'h0;
    if(slotValid) begin
      case(io_slot_opcode)
        4'b0010 : begin
          io_vectorWriteReqs_1_payload_addr = (io_slot_dest + 11'h001);
        end
        default : begin
        end
      endcase
    end
  end

  always @(*) begin
    io_vectorWriteReqs_1_payload_data = 32'h0;
    if(slotValid) begin
      case(io_slot_opcode)
        4'b0010 : begin
          io_vectorWriteReqs_1_payload_data = ((io_vCond_1 != 32'h0) ? io_vSrcA_1 : io_vSrcB_1);
        end
        default : begin
        end
      endcase
    end
  end

  always @(*) begin
    io_vectorWriteReqs_2_valid = 1'b0;
    if(slotValid) begin
      case(io_slot_opcode)
        4'b0010 : begin
          io_vectorWriteReqs_2_valid = 1'b1;
        end
        default : begin
        end
      endcase
    end
  end

  always @(*) begin
    io_vectorWriteReqs_2_payload_addr = 11'h0;
    if(slotValid) begin
      case(io_slot_opcode)
        4'b0010 : begin
          io_vectorWriteReqs_2_payload_addr = (io_slot_dest + 11'h002);
        end
        default : begin
        end
      endcase
    end
  end

  always @(*) begin
    io_vectorWriteReqs_2_payload_data = 32'h0;
    if(slotValid) begin
      case(io_slot_opcode)
        4'b0010 : begin
          io_vectorWriteReqs_2_payload_data = ((io_vCond_2 != 32'h0) ? io_vSrcA_2 : io_vSrcB_2);
        end
        default : begin
        end
      endcase
    end
  end

  always @(*) begin
    io_vectorWriteReqs_3_valid = 1'b0;
    if(slotValid) begin
      case(io_slot_opcode)
        4'b0010 : begin
          io_vectorWriteReqs_3_valid = 1'b1;
        end
        default : begin
        end
      endcase
    end
  end

  always @(*) begin
    io_vectorWriteReqs_3_payload_addr = 11'h0;
    if(slotValid) begin
      case(io_slot_opcode)
        4'b0010 : begin
          io_vectorWriteReqs_3_payload_addr = (io_slot_dest + 11'h003);
        end
        default : begin
        end
      endcase
    end
  end

  always @(*) begin
    io_vectorWriteReqs_3_payload_data = 32'h0;
    if(slotValid) begin
      case(io_slot_opcode)
        4'b0010 : begin
          io_vectorWriteReqs_3_payload_data = ((io_vCond_3 != 32'h0) ? io_vSrcA_3 : io_vSrcB_3);
        end
        default : begin
        end
      endcase
    end
  end

  always @(*) begin
    io_vectorWriteReqs_4_valid = 1'b0;
    if(slotValid) begin
      case(io_slot_opcode)
        4'b0010 : begin
          io_vectorWriteReqs_4_valid = 1'b1;
        end
        default : begin
        end
      endcase
    end
  end

  always @(*) begin
    io_vectorWriteReqs_4_payload_addr = 11'h0;
    if(slotValid) begin
      case(io_slot_opcode)
        4'b0010 : begin
          io_vectorWriteReqs_4_payload_addr = (io_slot_dest + 11'h004);
        end
        default : begin
        end
      endcase
    end
  end

  always @(*) begin
    io_vectorWriteReqs_4_payload_data = 32'h0;
    if(slotValid) begin
      case(io_slot_opcode)
        4'b0010 : begin
          io_vectorWriteReqs_4_payload_data = ((io_vCond_4 != 32'h0) ? io_vSrcA_4 : io_vSrcB_4);
        end
        default : begin
        end
      endcase
    end
  end

  always @(*) begin
    io_vectorWriteReqs_5_valid = 1'b0;
    if(slotValid) begin
      case(io_slot_opcode)
        4'b0010 : begin
          io_vectorWriteReqs_5_valid = 1'b1;
        end
        default : begin
        end
      endcase
    end
  end

  always @(*) begin
    io_vectorWriteReqs_5_payload_addr = 11'h0;
    if(slotValid) begin
      case(io_slot_opcode)
        4'b0010 : begin
          io_vectorWriteReqs_5_payload_addr = (io_slot_dest + 11'h005);
        end
        default : begin
        end
      endcase
    end
  end

  always @(*) begin
    io_vectorWriteReqs_5_payload_data = 32'h0;
    if(slotValid) begin
      case(io_slot_opcode)
        4'b0010 : begin
          io_vectorWriteReqs_5_payload_data = ((io_vCond_5 != 32'h0) ? io_vSrcA_5 : io_vSrcB_5);
        end
        default : begin
        end
      endcase
    end
  end

  always @(*) begin
    io_vectorWriteReqs_6_valid = 1'b0;
    if(slotValid) begin
      case(io_slot_opcode)
        4'b0010 : begin
          io_vectorWriteReqs_6_valid = 1'b1;
        end
        default : begin
        end
      endcase
    end
  end

  always @(*) begin
    io_vectorWriteReqs_6_payload_addr = 11'h0;
    if(slotValid) begin
      case(io_slot_opcode)
        4'b0010 : begin
          io_vectorWriteReqs_6_payload_addr = (io_slot_dest + 11'h006);
        end
        default : begin
        end
      endcase
    end
  end

  always @(*) begin
    io_vectorWriteReqs_6_payload_data = 32'h0;
    if(slotValid) begin
      case(io_slot_opcode)
        4'b0010 : begin
          io_vectorWriteReqs_6_payload_data = ((io_vCond_6 != 32'h0) ? io_vSrcA_6 : io_vSrcB_6);
        end
        default : begin
        end
      endcase
    end
  end

  always @(*) begin
    io_vectorWriteReqs_7_valid = 1'b0;
    if(slotValid) begin
      case(io_slot_opcode)
        4'b0010 : begin
          io_vectorWriteReqs_7_valid = 1'b1;
        end
        default : begin
        end
      endcase
    end
  end

  always @(*) begin
    io_vectorWriteReqs_7_payload_addr = 11'h0;
    if(slotValid) begin
      case(io_slot_opcode)
        4'b0010 : begin
          io_vectorWriteReqs_7_payload_addr = (io_slot_dest + 11'h007);
        end
        default : begin
        end
      endcase
    end
  end

  always @(*) begin
    io_vectorWriteReqs_7_payload_data = 32'h0;
    if(slotValid) begin
      case(io_slot_opcode)
        4'b0010 : begin
          io_vectorWriteReqs_7_payload_data = ((io_vCond_7 != 32'h0) ? io_vSrcA_7 : io_vSrcB_7);
        end
        default : begin
        end
      endcase
    end
  end

  always @(*) begin
    io_jumpTarget_valid = 1'b0;
    if(slotValid) begin
      case(io_slot_opcode)
        4'b0101 : begin
          if(when_FlowEngine_l109) begin
            io_jumpTarget_valid = 1'b1;
          end
        end
        4'b0110 : begin
          if(when_FlowEngine_l118) begin
            io_jumpTarget_valid = 1'b1;
          end
        end
        4'b0111 : begin
          io_jumpTarget_valid = 1'b1;
        end
        4'b1000 : begin
          io_jumpTarget_valid = 1'b1;
        end
        default : begin
        end
      endcase
    end
  end

  always @(*) begin
    io_jumpTarget_payload = 10'h0;
    if(slotValid) begin
      case(io_slot_opcode)
        4'b0101 : begin
          if(when_FlowEngine_l109) begin
            io_jumpTarget_payload = _zz_io_jumpTarget_payload[9:0];
          end
        end
        4'b0110 : begin
          if(when_FlowEngine_l118) begin
            io_jumpTarget_payload = _zz_io_jumpTarget_payload_1;
          end
        end
        4'b0111 : begin
          io_jumpTarget_payload = _zz_io_jumpTarget_payload_4[9:0];
        end
        4'b1000 : begin
          io_jumpTarget_payload = io_operandCond[9:0];
        end
        default : begin
        end
      endcase
    end
  end

  always @(*) begin
    io_halt = 1'b0;
    if(slotValid) begin
      case(io_slot_opcode)
        4'b0100 : begin
          io_halt = 1'b1;
        end
        default : begin
        end
      endcase
    end
  end

  assign when_FlowEngine_l109 = (io_operandCond != 32'h0);
  assign when_FlowEngine_l118 = (io_operandCond != 32'h0);

endmodule

module ValuEngine (
  input  wire          io_slots_0_valid,
  input  wire [3:0]    io_slots_0_opcode,
  input  wire [10:0]   io_slots_0_destBase,
  input  wire [10:0]   io_slots_0_src1Base,
  input  wire [10:0]   io_slots_0_src2Base,
  input  wire [10:0]   io_slots_0_src3Base,
  input  wire          io_valid,
  input  wire [31:0]   io_operandA_0_0,
  input  wire [31:0]   io_operandA_0_1,
  input  wire [31:0]   io_operandA_0_2,
  input  wire [31:0]   io_operandA_0_3,
  input  wire [31:0]   io_operandA_0_4,
  input  wire [31:0]   io_operandA_0_5,
  input  wire [31:0]   io_operandA_0_6,
  input  wire [31:0]   io_operandA_0_7,
  input  wire [31:0]   io_operandB_0_0,
  input  wire [31:0]   io_operandB_0_1,
  input  wire [31:0]   io_operandB_0_2,
  input  wire [31:0]   io_operandB_0_3,
  input  wire [31:0]   io_operandB_0_4,
  input  wire [31:0]   io_operandB_0_5,
  input  wire [31:0]   io_operandB_0_6,
  input  wire [31:0]   io_operandB_0_7,
  input  wire [31:0]   io_operandC_0_0,
  input  wire [31:0]   io_operandC_0_1,
  input  wire [31:0]   io_operandC_0_2,
  input  wire [31:0]   io_operandC_0_3,
  input  wire [31:0]   io_operandC_0_4,
  input  wire [31:0]   io_operandC_0_5,
  input  wire [31:0]   io_operandC_0_6,
  input  wire [31:0]   io_operandC_0_7,
  output wire          io_writeReqs_0_0_valid,
  output wire [10:0]   io_writeReqs_0_0_payload_addr,
  output wire [31:0]   io_writeReqs_0_0_payload_data,
  output wire          io_writeReqs_0_1_valid,
  output wire [10:0]   io_writeReqs_0_1_payload_addr,
  output wire [31:0]   io_writeReqs_0_1_payload_data,
  output wire          io_writeReqs_0_2_valid,
  output wire [10:0]   io_writeReqs_0_2_payload_addr,
  output wire [31:0]   io_writeReqs_0_2_payload_data,
  output wire          io_writeReqs_0_3_valid,
  output wire [10:0]   io_writeReqs_0_3_payload_addr,
  output wire [31:0]   io_writeReqs_0_3_payload_data,
  output wire          io_writeReqs_0_4_valid,
  output wire [10:0]   io_writeReqs_0_4_payload_addr,
  output wire [31:0]   io_writeReqs_0_4_payload_data,
  output wire          io_writeReqs_0_5_valid,
  output wire [10:0]   io_writeReqs_0_5_payload_addr,
  output wire [31:0]   io_writeReqs_0_5_payload_data,
  output wire          io_writeReqs_0_6_valid,
  output wire [10:0]   io_writeReqs_0_6_payload_addr,
  output wire [31:0]   io_writeReqs_0_6_payload_data,
  output wire          io_writeReqs_0_7_valid,
  output wire [10:0]   io_writeReqs_0_7_payload_addr,
  output wire [31:0]   io_writeReqs_0_7_payload_data,
  input  wire          clk,
  input  wire          reset
);

  wire                unsignedDivider_9_io_start;
  wire       [31:0]   unsignedDivider_9_io_dividend;
  wire                unsignedDivider_10_io_start;
  wire       [31:0]   unsignedDivider_10_io_dividend;
  wire                unsignedDivider_11_io_start;
  wire       [31:0]   unsignedDivider_11_io_dividend;
  wire                unsignedDivider_12_io_start;
  wire       [31:0]   unsignedDivider_12_io_dividend;
  wire                unsignedDivider_13_io_start;
  wire       [31:0]   unsignedDivider_13_io_dividend;
  wire                unsignedDivider_14_io_start;
  wire       [31:0]   unsignedDivider_14_io_dividend;
  wire                unsignedDivider_15_io_start;
  wire       [31:0]   unsignedDivider_15_io_dividend;
  wire                unsignedDivider_16_io_start;
  wire       [31:0]   unsignedDivider_16_io_dividend;
  wire                unsignedDivider_9_io_done;
  wire                unsignedDivider_9_io_busy;
  wire       [31:0]   unsignedDivider_9_io_quotient;
  wire       [31:0]   unsignedDivider_9_io_remainder;
  wire                unsignedDivider_10_io_done;
  wire                unsignedDivider_10_io_busy;
  wire       [31:0]   unsignedDivider_10_io_quotient;
  wire       [31:0]   unsignedDivider_10_io_remainder;
  wire                unsignedDivider_11_io_done;
  wire                unsignedDivider_11_io_busy;
  wire       [31:0]   unsignedDivider_11_io_quotient;
  wire       [31:0]   unsignedDivider_11_io_remainder;
  wire                unsignedDivider_12_io_done;
  wire                unsignedDivider_12_io_busy;
  wire       [31:0]   unsignedDivider_12_io_quotient;
  wire       [31:0]   unsignedDivider_12_io_remainder;
  wire                unsignedDivider_13_io_done;
  wire                unsignedDivider_13_io_busy;
  wire       [31:0]   unsignedDivider_13_io_quotient;
  wire       [31:0]   unsignedDivider_13_io_remainder;
  wire                unsignedDivider_14_io_done;
  wire                unsignedDivider_14_io_busy;
  wire       [31:0]   unsignedDivider_14_io_quotient;
  wire       [31:0]   unsignedDivider_14_io_remainder;
  wire                unsignedDivider_15_io_done;
  wire                unsignedDivider_15_io_busy;
  wire       [31:0]   unsignedDivider_15_io_quotient;
  wire       [31:0]   unsignedDivider_15_io_remainder;
  wire                unsignedDivider_16_io_done;
  wire                unsignedDivider_16_io_busy;
  wire       [31:0]   unsignedDivider_16_io_quotient;
  wire       [31:0]   unsignedDivider_16_io_remainder;
  wire       [31:0]   _zz_io_dividend;
  wire       [31:0]   _zz_io_dividend_1;
  wire       [63:0]   _zz__zz_io_writeReqs_0_0_payload_data_1;
  wire       [0:0]    _zz__zz_io_writeReqs_0_0_payload_data_1_1;
  wire       [0:0]    _zz__zz_io_writeReqs_0_0_payload_data_1_2;
  wire       [63:0]   _zz__zz_io_writeReqs_0_0_payload_data_1_3;
  wire       [63:0]   _zz__zz_io_writeReqs_0_0_payload_data_1_4;
  wire       [63:0]   _zz__zz_io_writeReqs_0_0_payload_data_1_5;
  wire       [10:0]   _zz_io_writeReqs_0_0_payload_addr_1;
  wire       [31:0]   _zz_io_dividend_2;
  wire       [31:0]   _zz_io_dividend_3;
  wire       [63:0]   _zz__zz_io_writeReqs_0_1_payload_data_1;
  wire       [0:0]    _zz__zz_io_writeReqs_0_1_payload_data_1_1;
  wire       [0:0]    _zz__zz_io_writeReqs_0_1_payload_data_1_2;
  wire       [63:0]   _zz__zz_io_writeReqs_0_1_payload_data_1_3;
  wire       [63:0]   _zz__zz_io_writeReqs_0_1_payload_data_1_4;
  wire       [63:0]   _zz__zz_io_writeReqs_0_1_payload_data_1_5;
  wire       [10:0]   _zz_io_writeReqs_0_1_payload_addr_1;
  wire       [31:0]   _zz_io_dividend_4;
  wire       [31:0]   _zz_io_dividend_5;
  wire       [63:0]   _zz__zz_io_writeReqs_0_2_payload_data_1;
  wire       [0:0]    _zz__zz_io_writeReqs_0_2_payload_data_1_1;
  wire       [0:0]    _zz__zz_io_writeReqs_0_2_payload_data_1_2;
  wire       [63:0]   _zz__zz_io_writeReqs_0_2_payload_data_1_3;
  wire       [63:0]   _zz__zz_io_writeReqs_0_2_payload_data_1_4;
  wire       [63:0]   _zz__zz_io_writeReqs_0_2_payload_data_1_5;
  wire       [10:0]   _zz_io_writeReqs_0_2_payload_addr_1;
  wire       [31:0]   _zz_io_dividend_6;
  wire       [31:0]   _zz_io_dividend_7;
  wire       [63:0]   _zz__zz_io_writeReqs_0_3_payload_data_1;
  wire       [0:0]    _zz__zz_io_writeReqs_0_3_payload_data_1_1;
  wire       [0:0]    _zz__zz_io_writeReqs_0_3_payload_data_1_2;
  wire       [63:0]   _zz__zz_io_writeReqs_0_3_payload_data_1_3;
  wire       [63:0]   _zz__zz_io_writeReqs_0_3_payload_data_1_4;
  wire       [63:0]   _zz__zz_io_writeReqs_0_3_payload_data_1_5;
  wire       [10:0]   _zz_io_writeReqs_0_3_payload_addr_1;
  wire       [31:0]   _zz_io_dividend_8;
  wire       [31:0]   _zz_io_dividend_9;
  wire       [63:0]   _zz__zz_io_writeReqs_0_4_payload_data_1;
  wire       [0:0]    _zz__zz_io_writeReqs_0_4_payload_data_1_1;
  wire       [0:0]    _zz__zz_io_writeReqs_0_4_payload_data_1_2;
  wire       [63:0]   _zz__zz_io_writeReqs_0_4_payload_data_1_3;
  wire       [63:0]   _zz__zz_io_writeReqs_0_4_payload_data_1_4;
  wire       [63:0]   _zz__zz_io_writeReqs_0_4_payload_data_1_5;
  wire       [10:0]   _zz_io_writeReqs_0_4_payload_addr_1;
  wire       [31:0]   _zz_io_dividend_10;
  wire       [31:0]   _zz_io_dividend_11;
  wire       [63:0]   _zz__zz_io_writeReqs_0_5_payload_data_1;
  wire       [0:0]    _zz__zz_io_writeReqs_0_5_payload_data_1_1;
  wire       [0:0]    _zz__zz_io_writeReqs_0_5_payload_data_1_2;
  wire       [63:0]   _zz__zz_io_writeReqs_0_5_payload_data_1_3;
  wire       [63:0]   _zz__zz_io_writeReqs_0_5_payload_data_1_4;
  wire       [63:0]   _zz__zz_io_writeReqs_0_5_payload_data_1_5;
  wire       [10:0]   _zz_io_writeReqs_0_5_payload_addr_1;
  wire       [31:0]   _zz_io_dividend_12;
  wire       [31:0]   _zz_io_dividend_13;
  wire       [63:0]   _zz__zz_io_writeReqs_0_6_payload_data_1;
  wire       [0:0]    _zz__zz_io_writeReqs_0_6_payload_data_1_1;
  wire       [0:0]    _zz__zz_io_writeReqs_0_6_payload_data_1_2;
  wire       [63:0]   _zz__zz_io_writeReqs_0_6_payload_data_1_3;
  wire       [63:0]   _zz__zz_io_writeReqs_0_6_payload_data_1_4;
  wire       [63:0]   _zz__zz_io_writeReqs_0_6_payload_data_1_5;
  wire       [10:0]   _zz_io_writeReqs_0_6_payload_addr_1;
  wire       [31:0]   _zz_io_dividend_14;
  wire       [31:0]   _zz_io_dividend_15;
  wire       [63:0]   _zz__zz_io_writeReqs_0_7_payload_data_1;
  wire       [0:0]    _zz__zz_io_writeReqs_0_7_payload_data_1_1;
  wire       [0:0]    _zz__zz_io_writeReqs_0_7_payload_data_1_2;
  wire       [63:0]   _zz__zz_io_writeReqs_0_7_payload_data_1_3;
  wire       [63:0]   _zz__zz_io_writeReqs_0_7_payload_data_1_4;
  wire       [63:0]   _zz__zz_io_writeReqs_0_7_payload_data_1_5;
  wire       [10:0]   _zz_io_writeReqs_0_7_payload_addr_1;
  wire                _zz_io_writeReqs_0_0_valid;
  reg        [10:0]   _zz_io_writeReqs_0_0_payload_addr;
  reg        [1:0]    _zz_io_writeReqs_0_0_payload_data;
  wire                _zz_io_writeReqs_0_0_valid_1;
  wire                when_ValuEngine_l72;
  wire                when_ValuEngine_l74;
  reg        [31:0]   _zz_io_writeReqs_0_0_payload_data_1;
  reg        [10:0]   _zz_io_writeReqs_0_1_payload_addr;
  reg        [1:0]    _zz_io_writeReqs_0_1_payload_data;
  wire                _zz_io_writeReqs_0_1_valid;
  wire                when_ValuEngine_l72_1;
  wire                when_ValuEngine_l74_1;
  reg        [31:0]   _zz_io_writeReqs_0_1_payload_data_1;
  reg        [10:0]   _zz_io_writeReqs_0_2_payload_addr;
  reg        [1:0]    _zz_io_writeReqs_0_2_payload_data;
  wire                _zz_io_writeReqs_0_2_valid;
  wire                when_ValuEngine_l72_2;
  wire                when_ValuEngine_l74_2;
  reg        [31:0]   _zz_io_writeReqs_0_2_payload_data_1;
  reg        [10:0]   _zz_io_writeReqs_0_3_payload_addr;
  reg        [1:0]    _zz_io_writeReqs_0_3_payload_data;
  wire                _zz_io_writeReqs_0_3_valid;
  wire                when_ValuEngine_l72_3;
  wire                when_ValuEngine_l74_3;
  reg        [31:0]   _zz_io_writeReqs_0_3_payload_data_1;
  reg        [10:0]   _zz_io_writeReqs_0_4_payload_addr;
  reg        [1:0]    _zz_io_writeReqs_0_4_payload_data;
  wire                _zz_io_writeReqs_0_4_valid;
  wire                when_ValuEngine_l72_4;
  wire                when_ValuEngine_l74_4;
  reg        [31:0]   _zz_io_writeReqs_0_4_payload_data_1;
  reg        [10:0]   _zz_io_writeReqs_0_5_payload_addr;
  reg        [1:0]    _zz_io_writeReqs_0_5_payload_data;
  wire                _zz_io_writeReqs_0_5_valid;
  wire                when_ValuEngine_l72_5;
  wire                when_ValuEngine_l74_5;
  reg        [31:0]   _zz_io_writeReqs_0_5_payload_data_1;
  reg        [10:0]   _zz_io_writeReqs_0_6_payload_addr;
  reg        [1:0]    _zz_io_writeReqs_0_6_payload_data;
  wire                _zz_io_writeReqs_0_6_valid;
  wire                when_ValuEngine_l72_6;
  wire                when_ValuEngine_l74_6;
  reg        [31:0]   _zz_io_writeReqs_0_6_payload_data_1;
  reg        [10:0]   _zz_io_writeReqs_0_7_payload_addr;
  reg        [1:0]    _zz_io_writeReqs_0_7_payload_data;
  wire                _zz_io_writeReqs_0_7_valid;
  wire                when_ValuEngine_l72_7;
  wire                when_ValuEngine_l74_7;
  reg        [31:0]   _zz_io_writeReqs_0_7_payload_data_1;

  assign _zz_io_dividend = (_zz_io_dividend_1 - 32'h00000001);
  assign _zz_io_dividend_1 = (io_operandA_0_0 + io_operandB_0_0);
  assign _zz__zz_io_writeReqs_0_0_payload_data_1 = (io_operandA_0_0 * io_operandB_0_0);
  assign _zz__zz_io_writeReqs_0_0_payload_data_1_1 = (io_operandA_0_0 < io_operandB_0_0);
  assign _zz__zz_io_writeReqs_0_0_payload_data_1_2 = (io_operandA_0_0 == io_operandB_0_0);
  assign _zz__zz_io_writeReqs_0_0_payload_data_1_3 = (_zz__zz_io_writeReqs_0_0_payload_data_1_4 + _zz__zz_io_writeReqs_0_0_payload_data_1_5);
  assign _zz__zz_io_writeReqs_0_0_payload_data_1_4 = (io_operandA_0_0 * io_operandB_0_0);
  assign _zz__zz_io_writeReqs_0_0_payload_data_1_5 = {32'd0, io_operandC_0_0};
  assign _zz_io_writeReqs_0_0_payload_addr_1 = (io_slots_0_destBase + 11'h0);
  assign _zz_io_dividend_2 = (_zz_io_dividend_3 - 32'h00000001);
  assign _zz_io_dividend_3 = (io_operandA_0_1 + io_operandB_0_1);
  assign _zz__zz_io_writeReqs_0_1_payload_data_1 = (io_operandA_0_1 * io_operandB_0_1);
  assign _zz__zz_io_writeReqs_0_1_payload_data_1_1 = (io_operandA_0_1 < io_operandB_0_1);
  assign _zz__zz_io_writeReqs_0_1_payload_data_1_2 = (io_operandA_0_1 == io_operandB_0_1);
  assign _zz__zz_io_writeReqs_0_1_payload_data_1_3 = (_zz__zz_io_writeReqs_0_1_payload_data_1_4 + _zz__zz_io_writeReqs_0_1_payload_data_1_5);
  assign _zz__zz_io_writeReqs_0_1_payload_data_1_4 = (io_operandA_0_1 * io_operandB_0_1);
  assign _zz__zz_io_writeReqs_0_1_payload_data_1_5 = {32'd0, io_operandC_0_1};
  assign _zz_io_writeReqs_0_1_payload_addr_1 = (io_slots_0_destBase + 11'h001);
  assign _zz_io_dividend_4 = (_zz_io_dividend_5 - 32'h00000001);
  assign _zz_io_dividend_5 = (io_operandA_0_2 + io_operandB_0_2);
  assign _zz__zz_io_writeReqs_0_2_payload_data_1 = (io_operandA_0_2 * io_operandB_0_2);
  assign _zz__zz_io_writeReqs_0_2_payload_data_1_1 = (io_operandA_0_2 < io_operandB_0_2);
  assign _zz__zz_io_writeReqs_0_2_payload_data_1_2 = (io_operandA_0_2 == io_operandB_0_2);
  assign _zz__zz_io_writeReqs_0_2_payload_data_1_3 = (_zz__zz_io_writeReqs_0_2_payload_data_1_4 + _zz__zz_io_writeReqs_0_2_payload_data_1_5);
  assign _zz__zz_io_writeReqs_0_2_payload_data_1_4 = (io_operandA_0_2 * io_operandB_0_2);
  assign _zz__zz_io_writeReqs_0_2_payload_data_1_5 = {32'd0, io_operandC_0_2};
  assign _zz_io_writeReqs_0_2_payload_addr_1 = (io_slots_0_destBase + 11'h002);
  assign _zz_io_dividend_6 = (_zz_io_dividend_7 - 32'h00000001);
  assign _zz_io_dividend_7 = (io_operandA_0_3 + io_operandB_0_3);
  assign _zz__zz_io_writeReqs_0_3_payload_data_1 = (io_operandA_0_3 * io_operandB_0_3);
  assign _zz__zz_io_writeReqs_0_3_payload_data_1_1 = (io_operandA_0_3 < io_operandB_0_3);
  assign _zz__zz_io_writeReqs_0_3_payload_data_1_2 = (io_operandA_0_3 == io_operandB_0_3);
  assign _zz__zz_io_writeReqs_0_3_payload_data_1_3 = (_zz__zz_io_writeReqs_0_3_payload_data_1_4 + _zz__zz_io_writeReqs_0_3_payload_data_1_5);
  assign _zz__zz_io_writeReqs_0_3_payload_data_1_4 = (io_operandA_0_3 * io_operandB_0_3);
  assign _zz__zz_io_writeReqs_0_3_payload_data_1_5 = {32'd0, io_operandC_0_3};
  assign _zz_io_writeReqs_0_3_payload_addr_1 = (io_slots_0_destBase + 11'h003);
  assign _zz_io_dividend_8 = (_zz_io_dividend_9 - 32'h00000001);
  assign _zz_io_dividend_9 = (io_operandA_0_4 + io_operandB_0_4);
  assign _zz__zz_io_writeReqs_0_4_payload_data_1 = (io_operandA_0_4 * io_operandB_0_4);
  assign _zz__zz_io_writeReqs_0_4_payload_data_1_1 = (io_operandA_0_4 < io_operandB_0_4);
  assign _zz__zz_io_writeReqs_0_4_payload_data_1_2 = (io_operandA_0_4 == io_operandB_0_4);
  assign _zz__zz_io_writeReqs_0_4_payload_data_1_3 = (_zz__zz_io_writeReqs_0_4_payload_data_1_4 + _zz__zz_io_writeReqs_0_4_payload_data_1_5);
  assign _zz__zz_io_writeReqs_0_4_payload_data_1_4 = (io_operandA_0_4 * io_operandB_0_4);
  assign _zz__zz_io_writeReqs_0_4_payload_data_1_5 = {32'd0, io_operandC_0_4};
  assign _zz_io_writeReqs_0_4_payload_addr_1 = (io_slots_0_destBase + 11'h004);
  assign _zz_io_dividend_10 = (_zz_io_dividend_11 - 32'h00000001);
  assign _zz_io_dividend_11 = (io_operandA_0_5 + io_operandB_0_5);
  assign _zz__zz_io_writeReqs_0_5_payload_data_1 = (io_operandA_0_5 * io_operandB_0_5);
  assign _zz__zz_io_writeReqs_0_5_payload_data_1_1 = (io_operandA_0_5 < io_operandB_0_5);
  assign _zz__zz_io_writeReqs_0_5_payload_data_1_2 = (io_operandA_0_5 == io_operandB_0_5);
  assign _zz__zz_io_writeReqs_0_5_payload_data_1_3 = (_zz__zz_io_writeReqs_0_5_payload_data_1_4 + _zz__zz_io_writeReqs_0_5_payload_data_1_5);
  assign _zz__zz_io_writeReqs_0_5_payload_data_1_4 = (io_operandA_0_5 * io_operandB_0_5);
  assign _zz__zz_io_writeReqs_0_5_payload_data_1_5 = {32'd0, io_operandC_0_5};
  assign _zz_io_writeReqs_0_5_payload_addr_1 = (io_slots_0_destBase + 11'h005);
  assign _zz_io_dividend_12 = (_zz_io_dividend_13 - 32'h00000001);
  assign _zz_io_dividend_13 = (io_operandA_0_6 + io_operandB_0_6);
  assign _zz__zz_io_writeReqs_0_6_payload_data_1 = (io_operandA_0_6 * io_operandB_0_6);
  assign _zz__zz_io_writeReqs_0_6_payload_data_1_1 = (io_operandA_0_6 < io_operandB_0_6);
  assign _zz__zz_io_writeReqs_0_6_payload_data_1_2 = (io_operandA_0_6 == io_operandB_0_6);
  assign _zz__zz_io_writeReqs_0_6_payload_data_1_3 = (_zz__zz_io_writeReqs_0_6_payload_data_1_4 + _zz__zz_io_writeReqs_0_6_payload_data_1_5);
  assign _zz__zz_io_writeReqs_0_6_payload_data_1_4 = (io_operandA_0_6 * io_operandB_0_6);
  assign _zz__zz_io_writeReqs_0_6_payload_data_1_5 = {32'd0, io_operandC_0_6};
  assign _zz_io_writeReqs_0_6_payload_addr_1 = (io_slots_0_destBase + 11'h006);
  assign _zz_io_dividend_14 = (_zz_io_dividend_15 - 32'h00000001);
  assign _zz_io_dividend_15 = (io_operandA_0_7 + io_operandB_0_7);
  assign _zz__zz_io_writeReqs_0_7_payload_data_1 = (io_operandA_0_7 * io_operandB_0_7);
  assign _zz__zz_io_writeReqs_0_7_payload_data_1_1 = (io_operandA_0_7 < io_operandB_0_7);
  assign _zz__zz_io_writeReqs_0_7_payload_data_1_2 = (io_operandA_0_7 == io_operandB_0_7);
  assign _zz__zz_io_writeReqs_0_7_payload_data_1_3 = (_zz__zz_io_writeReqs_0_7_payload_data_1_4 + _zz__zz_io_writeReqs_0_7_payload_data_1_5);
  assign _zz__zz_io_writeReqs_0_7_payload_data_1_4 = (io_operandA_0_7 * io_operandB_0_7);
  assign _zz__zz_io_writeReqs_0_7_payload_data_1_5 = {32'd0, io_operandC_0_7};
  assign _zz_io_writeReqs_0_7_payload_addr_1 = (io_slots_0_destBase + 11'h007);
  UnsignedDivider_8 unsignedDivider_9 (
    .io_start     (unsignedDivider_9_io_start          ), //i
    .io_dividend  (unsignedDivider_9_io_dividend[31:0] ), //i
    .io_divisor   (io_operandB_0_0[31:0]               ), //i
    .io_done      (unsignedDivider_9_io_done           ), //o
    .io_busy      (unsignedDivider_9_io_busy           ), //o
    .io_quotient  (unsignedDivider_9_io_quotient[31:0] ), //o
    .io_remainder (unsignedDivider_9_io_remainder[31:0]), //o
    .clk          (clk                                 ), //i
    .reset        (reset                               )  //i
  );
  UnsignedDivider_8 unsignedDivider_10 (
    .io_start     (unsignedDivider_10_io_start          ), //i
    .io_dividend  (unsignedDivider_10_io_dividend[31:0] ), //i
    .io_divisor   (io_operandB_0_1[31:0]                ), //i
    .io_done      (unsignedDivider_10_io_done           ), //o
    .io_busy      (unsignedDivider_10_io_busy           ), //o
    .io_quotient  (unsignedDivider_10_io_quotient[31:0] ), //o
    .io_remainder (unsignedDivider_10_io_remainder[31:0]), //o
    .clk          (clk                                  ), //i
    .reset        (reset                                )  //i
  );
  UnsignedDivider_8 unsignedDivider_11 (
    .io_start     (unsignedDivider_11_io_start          ), //i
    .io_dividend  (unsignedDivider_11_io_dividend[31:0] ), //i
    .io_divisor   (io_operandB_0_2[31:0]                ), //i
    .io_done      (unsignedDivider_11_io_done           ), //o
    .io_busy      (unsignedDivider_11_io_busy           ), //o
    .io_quotient  (unsignedDivider_11_io_quotient[31:0] ), //o
    .io_remainder (unsignedDivider_11_io_remainder[31:0]), //o
    .clk          (clk                                  ), //i
    .reset        (reset                                )  //i
  );
  UnsignedDivider_8 unsignedDivider_12 (
    .io_start     (unsignedDivider_12_io_start          ), //i
    .io_dividend  (unsignedDivider_12_io_dividend[31:0] ), //i
    .io_divisor   (io_operandB_0_3[31:0]                ), //i
    .io_done      (unsignedDivider_12_io_done           ), //o
    .io_busy      (unsignedDivider_12_io_busy           ), //o
    .io_quotient  (unsignedDivider_12_io_quotient[31:0] ), //o
    .io_remainder (unsignedDivider_12_io_remainder[31:0]), //o
    .clk          (clk                                  ), //i
    .reset        (reset                                )  //i
  );
  UnsignedDivider_8 unsignedDivider_13 (
    .io_start     (unsignedDivider_13_io_start          ), //i
    .io_dividend  (unsignedDivider_13_io_dividend[31:0] ), //i
    .io_divisor   (io_operandB_0_4[31:0]                ), //i
    .io_done      (unsignedDivider_13_io_done           ), //o
    .io_busy      (unsignedDivider_13_io_busy           ), //o
    .io_quotient  (unsignedDivider_13_io_quotient[31:0] ), //o
    .io_remainder (unsignedDivider_13_io_remainder[31:0]), //o
    .clk          (clk                                  ), //i
    .reset        (reset                                )  //i
  );
  UnsignedDivider_8 unsignedDivider_14 (
    .io_start     (unsignedDivider_14_io_start          ), //i
    .io_dividend  (unsignedDivider_14_io_dividend[31:0] ), //i
    .io_divisor   (io_operandB_0_5[31:0]                ), //i
    .io_done      (unsignedDivider_14_io_done           ), //o
    .io_busy      (unsignedDivider_14_io_busy           ), //o
    .io_quotient  (unsignedDivider_14_io_quotient[31:0] ), //o
    .io_remainder (unsignedDivider_14_io_remainder[31:0]), //o
    .clk          (clk                                  ), //i
    .reset        (reset                                )  //i
  );
  UnsignedDivider_8 unsignedDivider_15 (
    .io_start     (unsignedDivider_15_io_start          ), //i
    .io_dividend  (unsignedDivider_15_io_dividend[31:0] ), //i
    .io_divisor   (io_operandB_0_6[31:0]                ), //i
    .io_done      (unsignedDivider_15_io_done           ), //o
    .io_busy      (unsignedDivider_15_io_busy           ), //o
    .io_quotient  (unsignedDivider_15_io_quotient[31:0] ), //o
    .io_remainder (unsignedDivider_15_io_remainder[31:0]), //o
    .clk          (clk                                  ), //i
    .reset        (reset                                )  //i
  );
  UnsignedDivider_8 unsignedDivider_16 (
    .io_start     (unsignedDivider_16_io_start          ), //i
    .io_dividend  (unsignedDivider_16_io_dividend[31:0] ), //i
    .io_divisor   (io_operandB_0_7[31:0]                ), //i
    .io_done      (unsignedDivider_16_io_done           ), //o
    .io_busy      (unsignedDivider_16_io_busy           ), //o
    .io_quotient  (unsignedDivider_16_io_quotient[31:0] ), //o
    .io_remainder (unsignedDivider_16_io_remainder[31:0]), //o
    .clk          (clk                                  ), //i
    .reset        (reset                                )  //i
  );
  assign _zz_io_writeReqs_0_0_valid = (io_slots_0_valid && io_valid);
  assign _zz_io_writeReqs_0_0_valid_1 = (((io_slots_0_opcode == 4'b1010) || (io_slots_0_opcode == 4'b1011)) || (io_slots_0_opcode == 4'b1100));
  assign unsignedDivider_9_io_start = ((_zz_io_writeReqs_0_0_valid && _zz_io_writeReqs_0_0_valid_1) && (! unsignedDivider_9_io_busy));
  assign unsignedDivider_9_io_dividend = ((io_slots_0_opcode == 4'b1100) ? _zz_io_dividend : io_operandA_0_0);
  assign when_ValuEngine_l72 = (io_slots_0_opcode == 4'b1010);
  assign when_ValuEngine_l74 = (io_slots_0_opcode == 4'b1011);
  always @(*) begin
    _zz_io_writeReqs_0_0_payload_data_1 = 32'h0;
    case(io_slots_0_opcode)
      4'b0000 : begin
        _zz_io_writeReqs_0_0_payload_data_1 = (io_operandA_0_0 + io_operandB_0_0);
      end
      4'b0001 : begin
        _zz_io_writeReqs_0_0_payload_data_1 = (io_operandA_0_0 - io_operandB_0_0);
      end
      4'b0010 : begin
        _zz_io_writeReqs_0_0_payload_data_1 = _zz__zz_io_writeReqs_0_0_payload_data_1[31:0];
      end
      4'b0011 : begin
        _zz_io_writeReqs_0_0_payload_data_1 = (io_operandA_0_0 ^ io_operandB_0_0);
      end
      4'b0100 : begin
        _zz_io_writeReqs_0_0_payload_data_1 = (io_operandA_0_0 & io_operandB_0_0);
      end
      4'b0101 : begin
        _zz_io_writeReqs_0_0_payload_data_1 = (io_operandA_0_0 | io_operandB_0_0);
      end
      4'b0110 : begin
        _zz_io_writeReqs_0_0_payload_data_1 = (io_operandA_0_0 <<< io_operandB_0_0[4 : 0]);
      end
      4'b0111 : begin
        _zz_io_writeReqs_0_0_payload_data_1 = (io_operandA_0_0 >>> io_operandB_0_0[4 : 0]);
      end
      4'b1000 : begin
        _zz_io_writeReqs_0_0_payload_data_1 = {31'd0, _zz__zz_io_writeReqs_0_0_payload_data_1_1};
      end
      4'b1001 : begin
        _zz_io_writeReqs_0_0_payload_data_1 = {31'd0, _zz__zz_io_writeReqs_0_0_payload_data_1_2};
      end
      4'b1101 : begin
        _zz_io_writeReqs_0_0_payload_data_1 = io_operandC_0_0;
      end
      4'b1110 : begin
        _zz_io_writeReqs_0_0_payload_data_1 = _zz__zz_io_writeReqs_0_0_payload_data_1_3[31:0];
      end
      default : begin
      end
    endcase
  end

  assign io_writeReqs_0_0_valid = (unsignedDivider_9_io_done || (_zz_io_writeReqs_0_0_valid && (! _zz_io_writeReqs_0_0_valid_1)));
  assign io_writeReqs_0_0_payload_addr = (unsignedDivider_9_io_done ? _zz_io_writeReqs_0_0_payload_addr : _zz_io_writeReqs_0_0_payload_addr_1);
  assign io_writeReqs_0_0_payload_data = (unsignedDivider_9_io_done ? ((_zz_io_writeReqs_0_0_payload_data == 2'b00) ? unsignedDivider_9_io_remainder : unsignedDivider_9_io_quotient) : _zz_io_writeReqs_0_0_payload_data_1);
  assign _zz_io_writeReqs_0_1_valid = (((io_slots_0_opcode == 4'b1010) || (io_slots_0_opcode == 4'b1011)) || (io_slots_0_opcode == 4'b1100));
  assign unsignedDivider_10_io_start = ((_zz_io_writeReqs_0_0_valid && _zz_io_writeReqs_0_1_valid) && (! unsignedDivider_10_io_busy));
  assign unsignedDivider_10_io_dividend = ((io_slots_0_opcode == 4'b1100) ? _zz_io_dividend_2 : io_operandA_0_1);
  assign when_ValuEngine_l72_1 = (io_slots_0_opcode == 4'b1010);
  assign when_ValuEngine_l74_1 = (io_slots_0_opcode == 4'b1011);
  always @(*) begin
    _zz_io_writeReqs_0_1_payload_data_1 = 32'h0;
    case(io_slots_0_opcode)
      4'b0000 : begin
        _zz_io_writeReqs_0_1_payload_data_1 = (io_operandA_0_1 + io_operandB_0_1);
      end
      4'b0001 : begin
        _zz_io_writeReqs_0_1_payload_data_1 = (io_operandA_0_1 - io_operandB_0_1);
      end
      4'b0010 : begin
        _zz_io_writeReqs_0_1_payload_data_1 = _zz__zz_io_writeReqs_0_1_payload_data_1[31:0];
      end
      4'b0011 : begin
        _zz_io_writeReqs_0_1_payload_data_1 = (io_operandA_0_1 ^ io_operandB_0_1);
      end
      4'b0100 : begin
        _zz_io_writeReqs_0_1_payload_data_1 = (io_operandA_0_1 & io_operandB_0_1);
      end
      4'b0101 : begin
        _zz_io_writeReqs_0_1_payload_data_1 = (io_operandA_0_1 | io_operandB_0_1);
      end
      4'b0110 : begin
        _zz_io_writeReqs_0_1_payload_data_1 = (io_operandA_0_1 <<< io_operandB_0_1[4 : 0]);
      end
      4'b0111 : begin
        _zz_io_writeReqs_0_1_payload_data_1 = (io_operandA_0_1 >>> io_operandB_0_1[4 : 0]);
      end
      4'b1000 : begin
        _zz_io_writeReqs_0_1_payload_data_1 = {31'd0, _zz__zz_io_writeReqs_0_1_payload_data_1_1};
      end
      4'b1001 : begin
        _zz_io_writeReqs_0_1_payload_data_1 = {31'd0, _zz__zz_io_writeReqs_0_1_payload_data_1_2};
      end
      4'b1101 : begin
        _zz_io_writeReqs_0_1_payload_data_1 = io_operandC_0_0;
      end
      4'b1110 : begin
        _zz_io_writeReqs_0_1_payload_data_1 = _zz__zz_io_writeReqs_0_1_payload_data_1_3[31:0];
      end
      default : begin
      end
    endcase
  end

  assign io_writeReqs_0_1_valid = (unsignedDivider_10_io_done || (_zz_io_writeReqs_0_0_valid && (! _zz_io_writeReqs_0_1_valid)));
  assign io_writeReqs_0_1_payload_addr = (unsignedDivider_10_io_done ? _zz_io_writeReqs_0_1_payload_addr : _zz_io_writeReqs_0_1_payload_addr_1);
  assign io_writeReqs_0_1_payload_data = (unsignedDivider_10_io_done ? ((_zz_io_writeReqs_0_1_payload_data == 2'b00) ? unsignedDivider_10_io_remainder : unsignedDivider_10_io_quotient) : _zz_io_writeReqs_0_1_payload_data_1);
  assign _zz_io_writeReqs_0_2_valid = (((io_slots_0_opcode == 4'b1010) || (io_slots_0_opcode == 4'b1011)) || (io_slots_0_opcode == 4'b1100));
  assign unsignedDivider_11_io_start = ((_zz_io_writeReqs_0_0_valid && _zz_io_writeReqs_0_2_valid) && (! unsignedDivider_11_io_busy));
  assign unsignedDivider_11_io_dividend = ((io_slots_0_opcode == 4'b1100) ? _zz_io_dividend_4 : io_operandA_0_2);
  assign when_ValuEngine_l72_2 = (io_slots_0_opcode == 4'b1010);
  assign when_ValuEngine_l74_2 = (io_slots_0_opcode == 4'b1011);
  always @(*) begin
    _zz_io_writeReqs_0_2_payload_data_1 = 32'h0;
    case(io_slots_0_opcode)
      4'b0000 : begin
        _zz_io_writeReqs_0_2_payload_data_1 = (io_operandA_0_2 + io_operandB_0_2);
      end
      4'b0001 : begin
        _zz_io_writeReqs_0_2_payload_data_1 = (io_operandA_0_2 - io_operandB_0_2);
      end
      4'b0010 : begin
        _zz_io_writeReqs_0_2_payload_data_1 = _zz__zz_io_writeReqs_0_2_payload_data_1[31:0];
      end
      4'b0011 : begin
        _zz_io_writeReqs_0_2_payload_data_1 = (io_operandA_0_2 ^ io_operandB_0_2);
      end
      4'b0100 : begin
        _zz_io_writeReqs_0_2_payload_data_1 = (io_operandA_0_2 & io_operandB_0_2);
      end
      4'b0101 : begin
        _zz_io_writeReqs_0_2_payload_data_1 = (io_operandA_0_2 | io_operandB_0_2);
      end
      4'b0110 : begin
        _zz_io_writeReqs_0_2_payload_data_1 = (io_operandA_0_2 <<< io_operandB_0_2[4 : 0]);
      end
      4'b0111 : begin
        _zz_io_writeReqs_0_2_payload_data_1 = (io_operandA_0_2 >>> io_operandB_0_2[4 : 0]);
      end
      4'b1000 : begin
        _zz_io_writeReqs_0_2_payload_data_1 = {31'd0, _zz__zz_io_writeReqs_0_2_payload_data_1_1};
      end
      4'b1001 : begin
        _zz_io_writeReqs_0_2_payload_data_1 = {31'd0, _zz__zz_io_writeReqs_0_2_payload_data_1_2};
      end
      4'b1101 : begin
        _zz_io_writeReqs_0_2_payload_data_1 = io_operandC_0_0;
      end
      4'b1110 : begin
        _zz_io_writeReqs_0_2_payload_data_1 = _zz__zz_io_writeReqs_0_2_payload_data_1_3[31:0];
      end
      default : begin
      end
    endcase
  end

  assign io_writeReqs_0_2_valid = (unsignedDivider_11_io_done || (_zz_io_writeReqs_0_0_valid && (! _zz_io_writeReqs_0_2_valid)));
  assign io_writeReqs_0_2_payload_addr = (unsignedDivider_11_io_done ? _zz_io_writeReqs_0_2_payload_addr : _zz_io_writeReqs_0_2_payload_addr_1);
  assign io_writeReqs_0_2_payload_data = (unsignedDivider_11_io_done ? ((_zz_io_writeReqs_0_2_payload_data == 2'b00) ? unsignedDivider_11_io_remainder : unsignedDivider_11_io_quotient) : _zz_io_writeReqs_0_2_payload_data_1);
  assign _zz_io_writeReqs_0_3_valid = (((io_slots_0_opcode == 4'b1010) || (io_slots_0_opcode == 4'b1011)) || (io_slots_0_opcode == 4'b1100));
  assign unsignedDivider_12_io_start = ((_zz_io_writeReqs_0_0_valid && _zz_io_writeReqs_0_3_valid) && (! unsignedDivider_12_io_busy));
  assign unsignedDivider_12_io_dividend = ((io_slots_0_opcode == 4'b1100) ? _zz_io_dividend_6 : io_operandA_0_3);
  assign when_ValuEngine_l72_3 = (io_slots_0_opcode == 4'b1010);
  assign when_ValuEngine_l74_3 = (io_slots_0_opcode == 4'b1011);
  always @(*) begin
    _zz_io_writeReqs_0_3_payload_data_1 = 32'h0;
    case(io_slots_0_opcode)
      4'b0000 : begin
        _zz_io_writeReqs_0_3_payload_data_1 = (io_operandA_0_3 + io_operandB_0_3);
      end
      4'b0001 : begin
        _zz_io_writeReqs_0_3_payload_data_1 = (io_operandA_0_3 - io_operandB_0_3);
      end
      4'b0010 : begin
        _zz_io_writeReqs_0_3_payload_data_1 = _zz__zz_io_writeReqs_0_3_payload_data_1[31:0];
      end
      4'b0011 : begin
        _zz_io_writeReqs_0_3_payload_data_1 = (io_operandA_0_3 ^ io_operandB_0_3);
      end
      4'b0100 : begin
        _zz_io_writeReqs_0_3_payload_data_1 = (io_operandA_0_3 & io_operandB_0_3);
      end
      4'b0101 : begin
        _zz_io_writeReqs_0_3_payload_data_1 = (io_operandA_0_3 | io_operandB_0_3);
      end
      4'b0110 : begin
        _zz_io_writeReqs_0_3_payload_data_1 = (io_operandA_0_3 <<< io_operandB_0_3[4 : 0]);
      end
      4'b0111 : begin
        _zz_io_writeReqs_0_3_payload_data_1 = (io_operandA_0_3 >>> io_operandB_0_3[4 : 0]);
      end
      4'b1000 : begin
        _zz_io_writeReqs_0_3_payload_data_1 = {31'd0, _zz__zz_io_writeReqs_0_3_payload_data_1_1};
      end
      4'b1001 : begin
        _zz_io_writeReqs_0_3_payload_data_1 = {31'd0, _zz__zz_io_writeReqs_0_3_payload_data_1_2};
      end
      4'b1101 : begin
        _zz_io_writeReqs_0_3_payload_data_1 = io_operandC_0_0;
      end
      4'b1110 : begin
        _zz_io_writeReqs_0_3_payload_data_1 = _zz__zz_io_writeReqs_0_3_payload_data_1_3[31:0];
      end
      default : begin
      end
    endcase
  end

  assign io_writeReqs_0_3_valid = (unsignedDivider_12_io_done || (_zz_io_writeReqs_0_0_valid && (! _zz_io_writeReqs_0_3_valid)));
  assign io_writeReqs_0_3_payload_addr = (unsignedDivider_12_io_done ? _zz_io_writeReqs_0_3_payload_addr : _zz_io_writeReqs_0_3_payload_addr_1);
  assign io_writeReqs_0_3_payload_data = (unsignedDivider_12_io_done ? ((_zz_io_writeReqs_0_3_payload_data == 2'b00) ? unsignedDivider_12_io_remainder : unsignedDivider_12_io_quotient) : _zz_io_writeReqs_0_3_payload_data_1);
  assign _zz_io_writeReqs_0_4_valid = (((io_slots_0_opcode == 4'b1010) || (io_slots_0_opcode == 4'b1011)) || (io_slots_0_opcode == 4'b1100));
  assign unsignedDivider_13_io_start = ((_zz_io_writeReqs_0_0_valid && _zz_io_writeReqs_0_4_valid) && (! unsignedDivider_13_io_busy));
  assign unsignedDivider_13_io_dividend = ((io_slots_0_opcode == 4'b1100) ? _zz_io_dividend_8 : io_operandA_0_4);
  assign when_ValuEngine_l72_4 = (io_slots_0_opcode == 4'b1010);
  assign when_ValuEngine_l74_4 = (io_slots_0_opcode == 4'b1011);
  always @(*) begin
    _zz_io_writeReqs_0_4_payload_data_1 = 32'h0;
    case(io_slots_0_opcode)
      4'b0000 : begin
        _zz_io_writeReqs_0_4_payload_data_1 = (io_operandA_0_4 + io_operandB_0_4);
      end
      4'b0001 : begin
        _zz_io_writeReqs_0_4_payload_data_1 = (io_operandA_0_4 - io_operandB_0_4);
      end
      4'b0010 : begin
        _zz_io_writeReqs_0_4_payload_data_1 = _zz__zz_io_writeReqs_0_4_payload_data_1[31:0];
      end
      4'b0011 : begin
        _zz_io_writeReqs_0_4_payload_data_1 = (io_operandA_0_4 ^ io_operandB_0_4);
      end
      4'b0100 : begin
        _zz_io_writeReqs_0_4_payload_data_1 = (io_operandA_0_4 & io_operandB_0_4);
      end
      4'b0101 : begin
        _zz_io_writeReqs_0_4_payload_data_1 = (io_operandA_0_4 | io_operandB_0_4);
      end
      4'b0110 : begin
        _zz_io_writeReqs_0_4_payload_data_1 = (io_operandA_0_4 <<< io_operandB_0_4[4 : 0]);
      end
      4'b0111 : begin
        _zz_io_writeReqs_0_4_payload_data_1 = (io_operandA_0_4 >>> io_operandB_0_4[4 : 0]);
      end
      4'b1000 : begin
        _zz_io_writeReqs_0_4_payload_data_1 = {31'd0, _zz__zz_io_writeReqs_0_4_payload_data_1_1};
      end
      4'b1001 : begin
        _zz_io_writeReqs_0_4_payload_data_1 = {31'd0, _zz__zz_io_writeReqs_0_4_payload_data_1_2};
      end
      4'b1101 : begin
        _zz_io_writeReqs_0_4_payload_data_1 = io_operandC_0_0;
      end
      4'b1110 : begin
        _zz_io_writeReqs_0_4_payload_data_1 = _zz__zz_io_writeReqs_0_4_payload_data_1_3[31:0];
      end
      default : begin
      end
    endcase
  end

  assign io_writeReqs_0_4_valid = (unsignedDivider_13_io_done || (_zz_io_writeReqs_0_0_valid && (! _zz_io_writeReqs_0_4_valid)));
  assign io_writeReqs_0_4_payload_addr = (unsignedDivider_13_io_done ? _zz_io_writeReqs_0_4_payload_addr : _zz_io_writeReqs_0_4_payload_addr_1);
  assign io_writeReqs_0_4_payload_data = (unsignedDivider_13_io_done ? ((_zz_io_writeReqs_0_4_payload_data == 2'b00) ? unsignedDivider_13_io_remainder : unsignedDivider_13_io_quotient) : _zz_io_writeReqs_0_4_payload_data_1);
  assign _zz_io_writeReqs_0_5_valid = (((io_slots_0_opcode == 4'b1010) || (io_slots_0_opcode == 4'b1011)) || (io_slots_0_opcode == 4'b1100));
  assign unsignedDivider_14_io_start = ((_zz_io_writeReqs_0_0_valid && _zz_io_writeReqs_0_5_valid) && (! unsignedDivider_14_io_busy));
  assign unsignedDivider_14_io_dividend = ((io_slots_0_opcode == 4'b1100) ? _zz_io_dividend_10 : io_operandA_0_5);
  assign when_ValuEngine_l72_5 = (io_slots_0_opcode == 4'b1010);
  assign when_ValuEngine_l74_5 = (io_slots_0_opcode == 4'b1011);
  always @(*) begin
    _zz_io_writeReqs_0_5_payload_data_1 = 32'h0;
    case(io_slots_0_opcode)
      4'b0000 : begin
        _zz_io_writeReqs_0_5_payload_data_1 = (io_operandA_0_5 + io_operandB_0_5);
      end
      4'b0001 : begin
        _zz_io_writeReqs_0_5_payload_data_1 = (io_operandA_0_5 - io_operandB_0_5);
      end
      4'b0010 : begin
        _zz_io_writeReqs_0_5_payload_data_1 = _zz__zz_io_writeReqs_0_5_payload_data_1[31:0];
      end
      4'b0011 : begin
        _zz_io_writeReqs_0_5_payload_data_1 = (io_operandA_0_5 ^ io_operandB_0_5);
      end
      4'b0100 : begin
        _zz_io_writeReqs_0_5_payload_data_1 = (io_operandA_0_5 & io_operandB_0_5);
      end
      4'b0101 : begin
        _zz_io_writeReqs_0_5_payload_data_1 = (io_operandA_0_5 | io_operandB_0_5);
      end
      4'b0110 : begin
        _zz_io_writeReqs_0_5_payload_data_1 = (io_operandA_0_5 <<< io_operandB_0_5[4 : 0]);
      end
      4'b0111 : begin
        _zz_io_writeReqs_0_5_payload_data_1 = (io_operandA_0_5 >>> io_operandB_0_5[4 : 0]);
      end
      4'b1000 : begin
        _zz_io_writeReqs_0_5_payload_data_1 = {31'd0, _zz__zz_io_writeReqs_0_5_payload_data_1_1};
      end
      4'b1001 : begin
        _zz_io_writeReqs_0_5_payload_data_1 = {31'd0, _zz__zz_io_writeReqs_0_5_payload_data_1_2};
      end
      4'b1101 : begin
        _zz_io_writeReqs_0_5_payload_data_1 = io_operandC_0_0;
      end
      4'b1110 : begin
        _zz_io_writeReqs_0_5_payload_data_1 = _zz__zz_io_writeReqs_0_5_payload_data_1_3[31:0];
      end
      default : begin
      end
    endcase
  end

  assign io_writeReqs_0_5_valid = (unsignedDivider_14_io_done || (_zz_io_writeReqs_0_0_valid && (! _zz_io_writeReqs_0_5_valid)));
  assign io_writeReqs_0_5_payload_addr = (unsignedDivider_14_io_done ? _zz_io_writeReqs_0_5_payload_addr : _zz_io_writeReqs_0_5_payload_addr_1);
  assign io_writeReqs_0_5_payload_data = (unsignedDivider_14_io_done ? ((_zz_io_writeReqs_0_5_payload_data == 2'b00) ? unsignedDivider_14_io_remainder : unsignedDivider_14_io_quotient) : _zz_io_writeReqs_0_5_payload_data_1);
  assign _zz_io_writeReqs_0_6_valid = (((io_slots_0_opcode == 4'b1010) || (io_slots_0_opcode == 4'b1011)) || (io_slots_0_opcode == 4'b1100));
  assign unsignedDivider_15_io_start = ((_zz_io_writeReqs_0_0_valid && _zz_io_writeReqs_0_6_valid) && (! unsignedDivider_15_io_busy));
  assign unsignedDivider_15_io_dividend = ((io_slots_0_opcode == 4'b1100) ? _zz_io_dividend_12 : io_operandA_0_6);
  assign when_ValuEngine_l72_6 = (io_slots_0_opcode == 4'b1010);
  assign when_ValuEngine_l74_6 = (io_slots_0_opcode == 4'b1011);
  always @(*) begin
    _zz_io_writeReqs_0_6_payload_data_1 = 32'h0;
    case(io_slots_0_opcode)
      4'b0000 : begin
        _zz_io_writeReqs_0_6_payload_data_1 = (io_operandA_0_6 + io_operandB_0_6);
      end
      4'b0001 : begin
        _zz_io_writeReqs_0_6_payload_data_1 = (io_operandA_0_6 - io_operandB_0_6);
      end
      4'b0010 : begin
        _zz_io_writeReqs_0_6_payload_data_1 = _zz__zz_io_writeReqs_0_6_payload_data_1[31:0];
      end
      4'b0011 : begin
        _zz_io_writeReqs_0_6_payload_data_1 = (io_operandA_0_6 ^ io_operandB_0_6);
      end
      4'b0100 : begin
        _zz_io_writeReqs_0_6_payload_data_1 = (io_operandA_0_6 & io_operandB_0_6);
      end
      4'b0101 : begin
        _zz_io_writeReqs_0_6_payload_data_1 = (io_operandA_0_6 | io_operandB_0_6);
      end
      4'b0110 : begin
        _zz_io_writeReqs_0_6_payload_data_1 = (io_operandA_0_6 <<< io_operandB_0_6[4 : 0]);
      end
      4'b0111 : begin
        _zz_io_writeReqs_0_6_payload_data_1 = (io_operandA_0_6 >>> io_operandB_0_6[4 : 0]);
      end
      4'b1000 : begin
        _zz_io_writeReqs_0_6_payload_data_1 = {31'd0, _zz__zz_io_writeReqs_0_6_payload_data_1_1};
      end
      4'b1001 : begin
        _zz_io_writeReqs_0_6_payload_data_1 = {31'd0, _zz__zz_io_writeReqs_0_6_payload_data_1_2};
      end
      4'b1101 : begin
        _zz_io_writeReqs_0_6_payload_data_1 = io_operandC_0_0;
      end
      4'b1110 : begin
        _zz_io_writeReqs_0_6_payload_data_1 = _zz__zz_io_writeReqs_0_6_payload_data_1_3[31:0];
      end
      default : begin
      end
    endcase
  end

  assign io_writeReqs_0_6_valid = (unsignedDivider_15_io_done || (_zz_io_writeReqs_0_0_valid && (! _zz_io_writeReqs_0_6_valid)));
  assign io_writeReqs_0_6_payload_addr = (unsignedDivider_15_io_done ? _zz_io_writeReqs_0_6_payload_addr : _zz_io_writeReqs_0_6_payload_addr_1);
  assign io_writeReqs_0_6_payload_data = (unsignedDivider_15_io_done ? ((_zz_io_writeReqs_0_6_payload_data == 2'b00) ? unsignedDivider_15_io_remainder : unsignedDivider_15_io_quotient) : _zz_io_writeReqs_0_6_payload_data_1);
  assign _zz_io_writeReqs_0_7_valid = (((io_slots_0_opcode == 4'b1010) || (io_slots_0_opcode == 4'b1011)) || (io_slots_0_opcode == 4'b1100));
  assign unsignedDivider_16_io_start = ((_zz_io_writeReqs_0_0_valid && _zz_io_writeReqs_0_7_valid) && (! unsignedDivider_16_io_busy));
  assign unsignedDivider_16_io_dividend = ((io_slots_0_opcode == 4'b1100) ? _zz_io_dividend_14 : io_operandA_0_7);
  assign when_ValuEngine_l72_7 = (io_slots_0_opcode == 4'b1010);
  assign when_ValuEngine_l74_7 = (io_slots_0_opcode == 4'b1011);
  always @(*) begin
    _zz_io_writeReqs_0_7_payload_data_1 = 32'h0;
    case(io_slots_0_opcode)
      4'b0000 : begin
        _zz_io_writeReqs_0_7_payload_data_1 = (io_operandA_0_7 + io_operandB_0_7);
      end
      4'b0001 : begin
        _zz_io_writeReqs_0_7_payload_data_1 = (io_operandA_0_7 - io_operandB_0_7);
      end
      4'b0010 : begin
        _zz_io_writeReqs_0_7_payload_data_1 = _zz__zz_io_writeReqs_0_7_payload_data_1[31:0];
      end
      4'b0011 : begin
        _zz_io_writeReqs_0_7_payload_data_1 = (io_operandA_0_7 ^ io_operandB_0_7);
      end
      4'b0100 : begin
        _zz_io_writeReqs_0_7_payload_data_1 = (io_operandA_0_7 & io_operandB_0_7);
      end
      4'b0101 : begin
        _zz_io_writeReqs_0_7_payload_data_1 = (io_operandA_0_7 | io_operandB_0_7);
      end
      4'b0110 : begin
        _zz_io_writeReqs_0_7_payload_data_1 = (io_operandA_0_7 <<< io_operandB_0_7[4 : 0]);
      end
      4'b0111 : begin
        _zz_io_writeReqs_0_7_payload_data_1 = (io_operandA_0_7 >>> io_operandB_0_7[4 : 0]);
      end
      4'b1000 : begin
        _zz_io_writeReqs_0_7_payload_data_1 = {31'd0, _zz__zz_io_writeReqs_0_7_payload_data_1_1};
      end
      4'b1001 : begin
        _zz_io_writeReqs_0_7_payload_data_1 = {31'd0, _zz__zz_io_writeReqs_0_7_payload_data_1_2};
      end
      4'b1101 : begin
        _zz_io_writeReqs_0_7_payload_data_1 = io_operandC_0_0;
      end
      4'b1110 : begin
        _zz_io_writeReqs_0_7_payload_data_1 = _zz__zz_io_writeReqs_0_7_payload_data_1_3[31:0];
      end
      default : begin
      end
    endcase
  end

  assign io_writeReqs_0_7_valid = (unsignedDivider_16_io_done || (_zz_io_writeReqs_0_0_valid && (! _zz_io_writeReqs_0_7_valid)));
  assign io_writeReqs_0_7_payload_addr = (unsignedDivider_16_io_done ? _zz_io_writeReqs_0_7_payload_addr : _zz_io_writeReqs_0_7_payload_addr_1);
  assign io_writeReqs_0_7_payload_data = (unsignedDivider_16_io_done ? ((_zz_io_writeReqs_0_7_payload_data == 2'b00) ? unsignedDivider_16_io_remainder : unsignedDivider_16_io_quotient) : _zz_io_writeReqs_0_7_payload_data_1);
  always @(posedge clk) begin
    if(reset) begin
      _zz_io_writeReqs_0_0_payload_addr <= 11'h0;
      _zz_io_writeReqs_0_0_payload_data <= 2'b00;
      _zz_io_writeReqs_0_1_payload_addr <= 11'h0;
      _zz_io_writeReqs_0_1_payload_data <= 2'b00;
      _zz_io_writeReqs_0_2_payload_addr <= 11'h0;
      _zz_io_writeReqs_0_2_payload_data <= 2'b00;
      _zz_io_writeReqs_0_3_payload_addr <= 11'h0;
      _zz_io_writeReqs_0_3_payload_data <= 2'b00;
      _zz_io_writeReqs_0_4_payload_addr <= 11'h0;
      _zz_io_writeReqs_0_4_payload_data <= 2'b00;
      _zz_io_writeReqs_0_5_payload_addr <= 11'h0;
      _zz_io_writeReqs_0_5_payload_data <= 2'b00;
      _zz_io_writeReqs_0_6_payload_addr <= 11'h0;
      _zz_io_writeReqs_0_6_payload_data <= 2'b00;
      _zz_io_writeReqs_0_7_payload_addr <= 11'h0;
      _zz_io_writeReqs_0_7_payload_data <= 2'b00;
    end else begin
      if(unsignedDivider_9_io_start) begin
        _zz_io_writeReqs_0_0_payload_addr <= (io_slots_0_destBase + 11'h0);
        if(when_ValuEngine_l72) begin
          _zz_io_writeReqs_0_0_payload_data <= 2'b00;
        end else begin
          if(when_ValuEngine_l74) begin
            _zz_io_writeReqs_0_0_payload_data <= 2'b01;
          end else begin
            _zz_io_writeReqs_0_0_payload_data <= 2'b10;
          end
        end
      end
      if(unsignedDivider_10_io_start) begin
        _zz_io_writeReqs_0_1_payload_addr <= (io_slots_0_destBase + 11'h001);
        if(when_ValuEngine_l72_1) begin
          _zz_io_writeReqs_0_1_payload_data <= 2'b00;
        end else begin
          if(when_ValuEngine_l74_1) begin
            _zz_io_writeReqs_0_1_payload_data <= 2'b01;
          end else begin
            _zz_io_writeReqs_0_1_payload_data <= 2'b10;
          end
        end
      end
      if(unsignedDivider_11_io_start) begin
        _zz_io_writeReqs_0_2_payload_addr <= (io_slots_0_destBase + 11'h002);
        if(when_ValuEngine_l72_2) begin
          _zz_io_writeReqs_0_2_payload_data <= 2'b00;
        end else begin
          if(when_ValuEngine_l74_2) begin
            _zz_io_writeReqs_0_2_payload_data <= 2'b01;
          end else begin
            _zz_io_writeReqs_0_2_payload_data <= 2'b10;
          end
        end
      end
      if(unsignedDivider_12_io_start) begin
        _zz_io_writeReqs_0_3_payload_addr <= (io_slots_0_destBase + 11'h003);
        if(when_ValuEngine_l72_3) begin
          _zz_io_writeReqs_0_3_payload_data <= 2'b00;
        end else begin
          if(when_ValuEngine_l74_3) begin
            _zz_io_writeReqs_0_3_payload_data <= 2'b01;
          end else begin
            _zz_io_writeReqs_0_3_payload_data <= 2'b10;
          end
        end
      end
      if(unsignedDivider_13_io_start) begin
        _zz_io_writeReqs_0_4_payload_addr <= (io_slots_0_destBase + 11'h004);
        if(when_ValuEngine_l72_4) begin
          _zz_io_writeReqs_0_4_payload_data <= 2'b00;
        end else begin
          if(when_ValuEngine_l74_4) begin
            _zz_io_writeReqs_0_4_payload_data <= 2'b01;
          end else begin
            _zz_io_writeReqs_0_4_payload_data <= 2'b10;
          end
        end
      end
      if(unsignedDivider_14_io_start) begin
        _zz_io_writeReqs_0_5_payload_addr <= (io_slots_0_destBase + 11'h005);
        if(when_ValuEngine_l72_5) begin
          _zz_io_writeReqs_0_5_payload_data <= 2'b00;
        end else begin
          if(when_ValuEngine_l74_5) begin
            _zz_io_writeReqs_0_5_payload_data <= 2'b01;
          end else begin
            _zz_io_writeReqs_0_5_payload_data <= 2'b10;
          end
        end
      end
      if(unsignedDivider_15_io_start) begin
        _zz_io_writeReqs_0_6_payload_addr <= (io_slots_0_destBase + 11'h006);
        if(when_ValuEngine_l72_6) begin
          _zz_io_writeReqs_0_6_payload_data <= 2'b00;
        end else begin
          if(when_ValuEngine_l74_6) begin
            _zz_io_writeReqs_0_6_payload_data <= 2'b01;
          end else begin
            _zz_io_writeReqs_0_6_payload_data <= 2'b10;
          end
        end
      end
      if(unsignedDivider_16_io_start) begin
        _zz_io_writeReqs_0_7_payload_addr <= (io_slots_0_destBase + 11'h007);
        if(when_ValuEngine_l72_7) begin
          _zz_io_writeReqs_0_7_payload_data <= 2'b00;
        end else begin
          if(when_ValuEngine_l74_7) begin
            _zz_io_writeReqs_0_7_payload_data <= 2'b01;
          end else begin
            _zz_io_writeReqs_0_7_payload_data <= 2'b10;
          end
        end
      end
    end
  end


endmodule

module AluEngine (
  input  wire          io_slots_0_valid,
  input  wire [3:0]    io_slots_0_opcode,
  input  wire [10:0]   io_slots_0_dest,
  input  wire [10:0]   io_slots_0_src1,
  input  wire [10:0]   io_slots_0_src2,
  input  wire          io_valid,
  input  wire [31:0]   io_operandA_0,
  input  wire [31:0]   io_operandB_0,
  output wire          io_writeReqs_0_valid,
  output wire [10:0]   io_writeReqs_0_payload_addr,
  output wire [31:0]   io_writeReqs_0_payload_data,
  input  wire          clk,
  input  wire          reset
);

  wire                unsignedDivider_9_io_start;
  wire       [31:0]   unsignedDivider_9_io_dividend;
  wire                unsignedDivider_9_io_done;
  wire                unsignedDivider_9_io_busy;
  wire       [31:0]   unsignedDivider_9_io_quotient;
  wire       [31:0]   unsignedDivider_9_io_remainder;
  wire       [31:0]   _zz_io_dividend;
  wire       [31:0]   _zz_io_dividend_1;
  wire       [63:0]   _zz__zz_io_writeReqs_0_payload_data_1;
  wire       [0:0]    _zz__zz_io_writeReqs_0_payload_data_1_1;
  wire       [0:0]    _zz__zz_io_writeReqs_0_payload_data_1_2;
  wire                _zz_io_writeReqs_0_valid;
  reg        [10:0]   _zz_io_writeReqs_0_payload_addr;
  reg        [1:0]    _zz_io_writeReqs_0_payload_data;
  wire                _zz_io_writeReqs_0_valid_1;
  wire                when_AluEngine_l61;
  wire                when_AluEngine_l63;
  reg        [31:0]   _zz_io_writeReqs_0_payload_data_1;

  assign _zz_io_dividend = (_zz_io_dividend_1 - 32'h00000001);
  assign _zz_io_dividend_1 = (io_operandA_0 + io_operandB_0);
  assign _zz__zz_io_writeReqs_0_payload_data_1 = (io_operandA_0 * io_operandB_0);
  assign _zz__zz_io_writeReqs_0_payload_data_1_1 = (io_operandA_0 < io_operandB_0);
  assign _zz__zz_io_writeReqs_0_payload_data_1_2 = (io_operandA_0 == io_operandB_0);
  UnsignedDivider_8 unsignedDivider_9 (
    .io_start     (unsignedDivider_9_io_start          ), //i
    .io_dividend  (unsignedDivider_9_io_dividend[31:0] ), //i
    .io_divisor   (io_operandB_0[31:0]                 ), //i
    .io_done      (unsignedDivider_9_io_done           ), //o
    .io_busy      (unsignedDivider_9_io_busy           ), //o
    .io_quotient  (unsignedDivider_9_io_quotient[31:0] ), //o
    .io_remainder (unsignedDivider_9_io_remainder[31:0]), //o
    .clk          (clk                                 ), //i
    .reset        (reset                               )  //i
  );
  assign _zz_io_writeReqs_0_valid = (io_slots_0_valid && io_valid);
  assign _zz_io_writeReqs_0_valid_1 = (((io_slots_0_opcode == 4'b1010) || (io_slots_0_opcode == 4'b1011)) || (io_slots_0_opcode == 4'b1100));
  assign unsignedDivider_9_io_start = ((_zz_io_writeReqs_0_valid && _zz_io_writeReqs_0_valid_1) && (! unsignedDivider_9_io_busy));
  assign unsignedDivider_9_io_dividend = ((io_slots_0_opcode == 4'b1100) ? _zz_io_dividend : io_operandA_0);
  assign when_AluEngine_l61 = (io_slots_0_opcode == 4'b1010);
  assign when_AluEngine_l63 = (io_slots_0_opcode == 4'b1011);
  always @(*) begin
    _zz_io_writeReqs_0_payload_data_1 = 32'h0;
    case(io_slots_0_opcode)
      4'b0000 : begin
        _zz_io_writeReqs_0_payload_data_1 = (io_operandA_0 + io_operandB_0);
      end
      4'b0001 : begin
        _zz_io_writeReqs_0_payload_data_1 = (io_operandA_0 - io_operandB_0);
      end
      4'b0010 : begin
        _zz_io_writeReqs_0_payload_data_1 = _zz__zz_io_writeReqs_0_payload_data_1[31:0];
      end
      4'b0011 : begin
        _zz_io_writeReqs_0_payload_data_1 = (io_operandA_0 ^ io_operandB_0);
      end
      4'b0100 : begin
        _zz_io_writeReqs_0_payload_data_1 = (io_operandA_0 & io_operandB_0);
      end
      4'b0101 : begin
        _zz_io_writeReqs_0_payload_data_1 = (io_operandA_0 | io_operandB_0);
      end
      4'b0110 : begin
        _zz_io_writeReqs_0_payload_data_1 = (io_operandA_0 <<< io_operandB_0[4 : 0]);
      end
      4'b0111 : begin
        _zz_io_writeReqs_0_payload_data_1 = (io_operandA_0 >>> io_operandB_0[4 : 0]);
      end
      4'b1000 : begin
        _zz_io_writeReqs_0_payload_data_1 = {31'd0, _zz__zz_io_writeReqs_0_payload_data_1_1};
      end
      4'b1001 : begin
        _zz_io_writeReqs_0_payload_data_1 = {31'd0, _zz__zz_io_writeReqs_0_payload_data_1_2};
      end
      default : begin
      end
    endcase
  end

  assign io_writeReqs_0_valid = (unsignedDivider_9_io_done || (_zz_io_writeReqs_0_valid && (! _zz_io_writeReqs_0_valid_1)));
  assign io_writeReqs_0_payload_addr = (unsignedDivider_9_io_done ? _zz_io_writeReqs_0_payload_addr : io_slots_0_dest);
  assign io_writeReqs_0_payload_data = (unsignedDivider_9_io_done ? ((_zz_io_writeReqs_0_payload_data == 2'b00) ? unsignedDivider_9_io_remainder : unsignedDivider_9_io_quotient) : _zz_io_writeReqs_0_payload_data_1);
  always @(posedge clk) begin
    if(reset) begin
      _zz_io_writeReqs_0_payload_addr <= 11'h0;
      _zz_io_writeReqs_0_payload_data <= 2'b00;
    end else begin
      if(unsignedDivider_9_io_start) begin
        _zz_io_writeReqs_0_payload_addr <= io_slots_0_dest;
        if(when_AluEngine_l61) begin
          _zz_io_writeReqs_0_payload_data <= 2'b00;
        end else begin
          if(when_AluEngine_l63) begin
            _zz_io_writeReqs_0_payload_data <= 2'b01;
          end else begin
            _zz_io_writeReqs_0_payload_data <= 2'b10;
          end
        end
      end
    end
  end


endmodule

module BankedScratchMemory (
  input  wire [10:0]   io_valuReadAddr_0_0,
  input  wire [10:0]   io_valuReadAddr_0_1,
  input  wire [10:0]   io_valuReadAddr_0_2,
  input  wire [10:0]   io_valuReadAddr_0_3,
  input  wire [10:0]   io_valuReadAddr_0_4,
  input  wire [10:0]   io_valuReadAddr_0_5,
  input  wire [10:0]   io_valuReadAddr_0_6,
  input  wire [10:0]   io_valuReadAddr_0_7,
  input  wire [10:0]   io_valuReadAddr_1_0,
  input  wire [10:0]   io_valuReadAddr_1_1,
  input  wire [10:0]   io_valuReadAddr_1_2,
  input  wire [10:0]   io_valuReadAddr_1_3,
  input  wire [10:0]   io_valuReadAddr_1_4,
  input  wire [10:0]   io_valuReadAddr_1_5,
  input  wire [10:0]   io_valuReadAddr_1_6,
  input  wire [10:0]   io_valuReadAddr_1_7,
  input  wire          io_valuReadEn_0_0,
  input  wire          io_valuReadEn_0_1,
  input  wire          io_valuReadEn_0_2,
  input  wire          io_valuReadEn_0_3,
  input  wire          io_valuReadEn_0_4,
  input  wire          io_valuReadEn_0_5,
  input  wire          io_valuReadEn_0_6,
  input  wire          io_valuReadEn_0_7,
  input  wire          io_valuReadEn_1_0,
  input  wire          io_valuReadEn_1_1,
  input  wire          io_valuReadEn_1_2,
  input  wire          io_valuReadEn_1_3,
  input  wire          io_valuReadEn_1_4,
  input  wire          io_valuReadEn_1_5,
  input  wire          io_valuReadEn_1_6,
  input  wire          io_valuReadEn_1_7,
  output wire [31:0]   io_valuReadData_0_0,
  output wire [31:0]   io_valuReadData_0_1,
  output wire [31:0]   io_valuReadData_0_2,
  output wire [31:0]   io_valuReadData_0_3,
  output wire [31:0]   io_valuReadData_0_4,
  output wire [31:0]   io_valuReadData_0_5,
  output wire [31:0]   io_valuReadData_0_6,
  output wire [31:0]   io_valuReadData_0_7,
  output wire [31:0]   io_valuReadData_1_0,
  output wire [31:0]   io_valuReadData_1_1,
  output wire [31:0]   io_valuReadData_1_2,
  output wire [31:0]   io_valuReadData_1_3,
  output wire [31:0]   io_valuReadData_1_4,
  output wire [31:0]   io_valuReadData_1_5,
  output wire [31:0]   io_valuReadData_1_6,
  output wire [31:0]   io_valuReadData_1_7,
  input  wire [10:0]   io_scalarReadAddr_0,
  input  wire [10:0]   io_scalarReadAddr_1,
  input  wire [10:0]   io_scalarReadAddr_2,
  input  wire [10:0]   io_scalarReadAddr_3,
  input  wire [10:0]   io_scalarReadAddr_4,
  input  wire [10:0]   io_scalarReadAddr_5,
  input  wire [10:0]   io_scalarReadAddr_6,
  input  wire [10:0]   io_scalarReadAddr_7,
  input  wire [10:0]   io_scalarReadAddr_8,
  input  wire          io_scalarReadEn_0,
  input  wire          io_scalarReadEn_1,
  input  wire          io_scalarReadEn_2,
  input  wire          io_scalarReadEn_3,
  input  wire          io_scalarReadEn_4,
  input  wire          io_scalarReadEn_5,
  input  wire          io_scalarReadEn_6,
  input  wire          io_scalarReadEn_7,
  input  wire          io_scalarReadEn_8,
  output reg  [31:0]   io_scalarReadData_0,
  output reg  [31:0]   io_scalarReadData_1,
  output reg  [31:0]   io_scalarReadData_2,
  output reg  [31:0]   io_scalarReadData_3,
  output reg  [31:0]   io_scalarReadData_4,
  output reg  [31:0]   io_scalarReadData_5,
  output reg  [31:0]   io_scalarReadData_6,
  output reg  [31:0]   io_scalarReadData_7,
  output reg  [31:0]   io_scalarReadData_8,
  input  wire [10:0]   io_writeAddr_0,
  input  wire [10:0]   io_writeAddr_1,
  input  wire [10:0]   io_writeAddr_2,
  input  wire [10:0]   io_writeAddr_3,
  input  wire [10:0]   io_writeAddr_4,
  input  wire [10:0]   io_writeAddr_5,
  input  wire [10:0]   io_writeAddr_6,
  input  wire [10:0]   io_writeAddr_7,
  input  wire [10:0]   io_writeAddr_8,
  input  wire [10:0]   io_writeAddr_9,
  input  wire [10:0]   io_writeAddr_10,
  input  wire [10:0]   io_writeAddr_11,
  input  wire [10:0]   io_writeAddr_12,
  input  wire [10:0]   io_writeAddr_13,
  input  wire [10:0]   io_writeAddr_14,
  input  wire [10:0]   io_writeAddr_15,
  input  wire [10:0]   io_writeAddr_16,
  input  wire [10:0]   io_writeAddr_17,
  input  wire [10:0]   io_writeAddr_18,
  input  wire [10:0]   io_writeAddr_19,
  input  wire [10:0]   io_writeAddr_20,
  input  wire [10:0]   io_writeAddr_21,
  input  wire [10:0]   io_writeAddr_22,
  input  wire [10:0]   io_writeAddr_23,
  input  wire [10:0]   io_writeAddr_24,
  input  wire [10:0]   io_writeAddr_25,
  input  wire [10:0]   io_writeAddr_26,
  input  wire [10:0]   io_writeAddr_27,
  input  wire [31:0]   io_writeData_0,
  input  wire [31:0]   io_writeData_1,
  input  wire [31:0]   io_writeData_2,
  input  wire [31:0]   io_writeData_3,
  input  wire [31:0]   io_writeData_4,
  input  wire [31:0]   io_writeData_5,
  input  wire [31:0]   io_writeData_6,
  input  wire [31:0]   io_writeData_7,
  input  wire [31:0]   io_writeData_8,
  input  wire [31:0]   io_writeData_9,
  input  wire [31:0]   io_writeData_10,
  input  wire [31:0]   io_writeData_11,
  input  wire [31:0]   io_writeData_12,
  input  wire [31:0]   io_writeData_13,
  input  wire [31:0]   io_writeData_14,
  input  wire [31:0]   io_writeData_15,
  input  wire [31:0]   io_writeData_16,
  input  wire [31:0]   io_writeData_17,
  input  wire [31:0]   io_writeData_18,
  input  wire [31:0]   io_writeData_19,
  input  wire [31:0]   io_writeData_20,
  input  wire [31:0]   io_writeData_21,
  input  wire [31:0]   io_writeData_22,
  input  wire [31:0]   io_writeData_23,
  input  wire [31:0]   io_writeData_24,
  input  wire [31:0]   io_writeData_25,
  input  wire [31:0]   io_writeData_26,
  input  wire [31:0]   io_writeData_27,
  input  wire          io_writeEn_0,
  input  wire          io_writeEn_1,
  input  wire          io_writeEn_2,
  input  wire          io_writeEn_3,
  input  wire          io_writeEn_4,
  input  wire          io_writeEn_5,
  input  wire          io_writeEn_6,
  input  wire          io_writeEn_7,
  input  wire          io_writeEn_8,
  input  wire          io_writeEn_9,
  input  wire          io_writeEn_10,
  input  wire          io_writeEn_11,
  input  wire          io_writeEn_12,
  input  wire          io_writeEn_13,
  input  wire          io_writeEn_14,
  input  wire          io_writeEn_15,
  input  wire          io_writeEn_16,
  input  wire          io_writeEn_17,
  input  wire          io_writeEn_18,
  input  wire          io_writeEn_19,
  input  wire          io_writeEn_20,
  input  wire          io_writeEn_21,
  input  wire          io_writeEn_22,
  input  wire          io_writeEn_23,
  input  wire          io_writeEn_24,
  input  wire          io_writeEn_25,
  input  wire          io_writeEn_26,
  input  wire          io_writeEn_27,
  output reg           io_conflict,
  input  wire          clk,
  input  wire          reset
);

  reg        [7:0]    banks_0_io_reads_0_addr;
  reg                 banks_0_io_reads_0_en;
  reg        [7:0]    banks_0_io_reads_1_addr;
  reg                 banks_0_io_reads_1_en;
  reg        [7:0]    banks_0_io_reads_2_addr;
  reg                 banks_0_io_reads_2_en;
  reg        [7:0]    banks_0_io_write_addr;
  reg        [31:0]   banks_0_io_write_data;
  reg                 banks_0_io_write_en;
  reg        [7:0]    banks_1_io_reads_0_addr;
  reg                 banks_1_io_reads_0_en;
  reg        [7:0]    banks_1_io_reads_1_addr;
  reg                 banks_1_io_reads_1_en;
  reg        [7:0]    banks_1_io_reads_2_addr;
  reg                 banks_1_io_reads_2_en;
  reg        [7:0]    banks_1_io_write_addr;
  reg        [31:0]   banks_1_io_write_data;
  reg                 banks_1_io_write_en;
  reg        [7:0]    banks_2_io_reads_0_addr;
  reg                 banks_2_io_reads_0_en;
  reg        [7:0]    banks_2_io_reads_1_addr;
  reg                 banks_2_io_reads_1_en;
  reg        [7:0]    banks_2_io_reads_2_addr;
  reg                 banks_2_io_reads_2_en;
  reg        [7:0]    banks_2_io_write_addr;
  reg        [31:0]   banks_2_io_write_data;
  reg                 banks_2_io_write_en;
  reg        [7:0]    banks_3_io_reads_0_addr;
  reg                 banks_3_io_reads_0_en;
  reg        [7:0]    banks_3_io_reads_1_addr;
  reg                 banks_3_io_reads_1_en;
  reg        [7:0]    banks_3_io_reads_2_addr;
  reg                 banks_3_io_reads_2_en;
  reg        [7:0]    banks_3_io_write_addr;
  reg        [31:0]   banks_3_io_write_data;
  reg                 banks_3_io_write_en;
  reg        [7:0]    banks_4_io_reads_0_addr;
  reg                 banks_4_io_reads_0_en;
  reg        [7:0]    banks_4_io_reads_1_addr;
  reg                 banks_4_io_reads_1_en;
  reg        [7:0]    banks_4_io_reads_2_addr;
  reg                 banks_4_io_reads_2_en;
  reg        [7:0]    banks_4_io_write_addr;
  reg        [31:0]   banks_4_io_write_data;
  reg                 banks_4_io_write_en;
  reg        [7:0]    banks_5_io_reads_0_addr;
  reg                 banks_5_io_reads_0_en;
  reg        [7:0]    banks_5_io_reads_1_addr;
  reg                 banks_5_io_reads_1_en;
  reg        [7:0]    banks_5_io_reads_2_addr;
  reg                 banks_5_io_reads_2_en;
  reg        [7:0]    banks_5_io_write_addr;
  reg        [31:0]   banks_5_io_write_data;
  reg                 banks_5_io_write_en;
  reg        [7:0]    banks_6_io_reads_0_addr;
  reg                 banks_6_io_reads_0_en;
  reg        [7:0]    banks_6_io_reads_1_addr;
  reg                 banks_6_io_reads_1_en;
  reg        [7:0]    banks_6_io_reads_2_addr;
  reg                 banks_6_io_reads_2_en;
  reg        [7:0]    banks_6_io_write_addr;
  reg        [31:0]   banks_6_io_write_data;
  reg                 banks_6_io_write_en;
  reg        [7:0]    banks_7_io_reads_0_addr;
  reg                 banks_7_io_reads_0_en;
  reg        [7:0]    banks_7_io_reads_1_addr;
  reg                 banks_7_io_reads_1_en;
  reg        [7:0]    banks_7_io_reads_2_addr;
  reg                 banks_7_io_reads_2_en;
  reg        [7:0]    banks_7_io_write_addr;
  reg        [31:0]   banks_7_io_write_data;
  reg                 banks_7_io_write_en;
  wire       [31:0]   banks_0_io_reads_0_data;
  wire       [31:0]   banks_0_io_reads_1_data;
  wire       [31:0]   banks_0_io_reads_2_data;
  wire       [31:0]   banks_1_io_reads_0_data;
  wire       [31:0]   banks_1_io_reads_1_data;
  wire       [31:0]   banks_1_io_reads_2_data;
  wire       [31:0]   banks_2_io_reads_0_data;
  wire       [31:0]   banks_2_io_reads_1_data;
  wire       [31:0]   banks_2_io_reads_2_data;
  wire       [31:0]   banks_3_io_reads_0_data;
  wire       [31:0]   banks_3_io_reads_1_data;
  wire       [31:0]   banks_3_io_reads_2_data;
  wire       [31:0]   banks_4_io_reads_0_data;
  wire       [31:0]   banks_4_io_reads_1_data;
  wire       [31:0]   banks_4_io_reads_2_data;
  wire       [31:0]   banks_5_io_reads_0_data;
  wire       [31:0]   banks_5_io_reads_1_data;
  wire       [31:0]   banks_5_io_reads_2_data;
  wire       [31:0]   banks_6_io_reads_0_data;
  wire       [31:0]   banks_6_io_reads_1_data;
  wire       [31:0]   banks_6_io_reads_2_data;
  wire       [31:0]   banks_7_io_reads_0_data;
  wire       [31:0]   banks_7_io_reads_1_data;
  wire       [31:0]   banks_7_io_reads_2_data;
  wire                _zz__zz_when_BankedScratchMemory_l203_7;
  wire                _zz__zz_when_BankedScratchMemory_l203_7_1;
  wire                _zz__zz_when_BankedScratchMemory_l203_8;
  wire                _zz__zz_when_BankedScratchMemory_l203_8_1;
  wire                _zz__zz_when_BankedScratchMemory_l203_8_2;
  wire       [2:0]    _zz_when_BankedScratchMemory_l160;
  wire       [7:0]    _zz_io_reads_0_addr;
  reg        [31:0]   _zz_io_valuReadData_0_0;
  wire                when_BankedScratchMemory_l160;
  wire                when_BankedScratchMemory_l160_1;
  wire                when_BankedScratchMemory_l160_2;
  wire                when_BankedScratchMemory_l160_3;
  wire                when_BankedScratchMemory_l160_4;
  wire                when_BankedScratchMemory_l160_5;
  wire                when_BankedScratchMemory_l160_6;
  wire                when_BankedScratchMemory_l160_7;
  wire       [2:0]    _zz_when_BankedScratchMemory_l160_1;
  wire       [7:0]    _zz_io_reads_0_addr_1;
  reg        [31:0]   _zz_io_valuReadData_0_1;
  wire                when_BankedScratchMemory_l160_8;
  wire                when_BankedScratchMemory_l160_9;
  wire                when_BankedScratchMemory_l160_10;
  wire                when_BankedScratchMemory_l160_11;
  wire                when_BankedScratchMemory_l160_12;
  wire                when_BankedScratchMemory_l160_13;
  wire                when_BankedScratchMemory_l160_14;
  wire                when_BankedScratchMemory_l160_15;
  wire       [2:0]    _zz_when_BankedScratchMemory_l160_2;
  wire       [7:0]    _zz_io_reads_0_addr_2;
  reg        [31:0]   _zz_io_valuReadData_0_2;
  wire                when_BankedScratchMemory_l160_16;
  wire                when_BankedScratchMemory_l160_17;
  wire                when_BankedScratchMemory_l160_18;
  wire                when_BankedScratchMemory_l160_19;
  wire                when_BankedScratchMemory_l160_20;
  wire                when_BankedScratchMemory_l160_21;
  wire                when_BankedScratchMemory_l160_22;
  wire                when_BankedScratchMemory_l160_23;
  wire       [2:0]    _zz_when_BankedScratchMemory_l160_3;
  wire       [7:0]    _zz_io_reads_0_addr_3;
  reg        [31:0]   _zz_io_valuReadData_0_3;
  wire                when_BankedScratchMemory_l160_24;
  wire                when_BankedScratchMemory_l160_25;
  wire                when_BankedScratchMemory_l160_26;
  wire                when_BankedScratchMemory_l160_27;
  wire                when_BankedScratchMemory_l160_28;
  wire                when_BankedScratchMemory_l160_29;
  wire                when_BankedScratchMemory_l160_30;
  wire                when_BankedScratchMemory_l160_31;
  wire       [2:0]    _zz_when_BankedScratchMemory_l160_4;
  wire       [7:0]    _zz_io_reads_0_addr_4;
  reg        [31:0]   _zz_io_valuReadData_0_4;
  wire                when_BankedScratchMemory_l160_32;
  wire                when_BankedScratchMemory_l160_33;
  wire                when_BankedScratchMemory_l160_34;
  wire                when_BankedScratchMemory_l160_35;
  wire                when_BankedScratchMemory_l160_36;
  wire                when_BankedScratchMemory_l160_37;
  wire                when_BankedScratchMemory_l160_38;
  wire                when_BankedScratchMemory_l160_39;
  wire       [2:0]    _zz_when_BankedScratchMemory_l160_5;
  wire       [7:0]    _zz_io_reads_0_addr_5;
  reg        [31:0]   _zz_io_valuReadData_0_5;
  wire                when_BankedScratchMemory_l160_40;
  wire                when_BankedScratchMemory_l160_41;
  wire                when_BankedScratchMemory_l160_42;
  wire                when_BankedScratchMemory_l160_43;
  wire                when_BankedScratchMemory_l160_44;
  wire                when_BankedScratchMemory_l160_45;
  wire                when_BankedScratchMemory_l160_46;
  wire                when_BankedScratchMemory_l160_47;
  wire       [2:0]    _zz_when_BankedScratchMemory_l160_6;
  wire       [7:0]    _zz_io_reads_0_addr_6;
  reg        [31:0]   _zz_io_valuReadData_0_6;
  wire                when_BankedScratchMemory_l160_48;
  wire                when_BankedScratchMemory_l160_49;
  wire                when_BankedScratchMemory_l160_50;
  wire                when_BankedScratchMemory_l160_51;
  wire                when_BankedScratchMemory_l160_52;
  wire                when_BankedScratchMemory_l160_53;
  wire                when_BankedScratchMemory_l160_54;
  wire                when_BankedScratchMemory_l160_55;
  wire       [2:0]    _zz_when_BankedScratchMemory_l160_7;
  wire       [7:0]    _zz_io_reads_0_addr_7;
  reg        [31:0]   _zz_io_valuReadData_0_7;
  wire                when_BankedScratchMemory_l160_56;
  wire                when_BankedScratchMemory_l160_57;
  wire                when_BankedScratchMemory_l160_58;
  wire                when_BankedScratchMemory_l160_59;
  wire                when_BankedScratchMemory_l160_60;
  wire                when_BankedScratchMemory_l160_61;
  wire                when_BankedScratchMemory_l160_62;
  wire                when_BankedScratchMemory_l160_63;
  wire       [2:0]    _zz_when_BankedScratchMemory_l160_8;
  wire       [7:0]    _zz_io_reads_1_addr;
  reg        [31:0]   _zz_io_valuReadData_1_0;
  wire                when_BankedScratchMemory_l160_64;
  wire                when_BankedScratchMemory_l160_65;
  wire                when_BankedScratchMemory_l160_66;
  wire                when_BankedScratchMemory_l160_67;
  wire                when_BankedScratchMemory_l160_68;
  wire                when_BankedScratchMemory_l160_69;
  wire                when_BankedScratchMemory_l160_70;
  wire                when_BankedScratchMemory_l160_71;
  wire       [2:0]    _zz_when_BankedScratchMemory_l160_9;
  wire       [7:0]    _zz_io_reads_1_addr_1;
  reg        [31:0]   _zz_io_valuReadData_1_1;
  wire                when_BankedScratchMemory_l160_72;
  wire                when_BankedScratchMemory_l160_73;
  wire                when_BankedScratchMemory_l160_74;
  wire                when_BankedScratchMemory_l160_75;
  wire                when_BankedScratchMemory_l160_76;
  wire                when_BankedScratchMemory_l160_77;
  wire                when_BankedScratchMemory_l160_78;
  wire                when_BankedScratchMemory_l160_79;
  wire       [2:0]    _zz_when_BankedScratchMemory_l160_10;
  wire       [7:0]    _zz_io_reads_1_addr_2;
  reg        [31:0]   _zz_io_valuReadData_1_2;
  wire                when_BankedScratchMemory_l160_80;
  wire                when_BankedScratchMemory_l160_81;
  wire                when_BankedScratchMemory_l160_82;
  wire                when_BankedScratchMemory_l160_83;
  wire                when_BankedScratchMemory_l160_84;
  wire                when_BankedScratchMemory_l160_85;
  wire                when_BankedScratchMemory_l160_86;
  wire                when_BankedScratchMemory_l160_87;
  wire       [2:0]    _zz_when_BankedScratchMemory_l160_11;
  wire       [7:0]    _zz_io_reads_1_addr_3;
  reg        [31:0]   _zz_io_valuReadData_1_3;
  wire                when_BankedScratchMemory_l160_88;
  wire                when_BankedScratchMemory_l160_89;
  wire                when_BankedScratchMemory_l160_90;
  wire                when_BankedScratchMemory_l160_91;
  wire                when_BankedScratchMemory_l160_92;
  wire                when_BankedScratchMemory_l160_93;
  wire                when_BankedScratchMemory_l160_94;
  wire                when_BankedScratchMemory_l160_95;
  wire       [2:0]    _zz_when_BankedScratchMemory_l160_12;
  wire       [7:0]    _zz_io_reads_1_addr_4;
  reg        [31:0]   _zz_io_valuReadData_1_4;
  wire                when_BankedScratchMemory_l160_96;
  wire                when_BankedScratchMemory_l160_97;
  wire                when_BankedScratchMemory_l160_98;
  wire                when_BankedScratchMemory_l160_99;
  wire                when_BankedScratchMemory_l160_100;
  wire                when_BankedScratchMemory_l160_101;
  wire                when_BankedScratchMemory_l160_102;
  wire                when_BankedScratchMemory_l160_103;
  wire       [2:0]    _zz_when_BankedScratchMemory_l160_13;
  wire       [7:0]    _zz_io_reads_1_addr_5;
  reg        [31:0]   _zz_io_valuReadData_1_5;
  wire                when_BankedScratchMemory_l160_104;
  wire                when_BankedScratchMemory_l160_105;
  wire                when_BankedScratchMemory_l160_106;
  wire                when_BankedScratchMemory_l160_107;
  wire                when_BankedScratchMemory_l160_108;
  wire                when_BankedScratchMemory_l160_109;
  wire                when_BankedScratchMemory_l160_110;
  wire                when_BankedScratchMemory_l160_111;
  wire       [2:0]    _zz_when_BankedScratchMemory_l160_14;
  wire       [7:0]    _zz_io_reads_1_addr_6;
  reg        [31:0]   _zz_io_valuReadData_1_6;
  wire                when_BankedScratchMemory_l160_112;
  wire                when_BankedScratchMemory_l160_113;
  wire                when_BankedScratchMemory_l160_114;
  wire                when_BankedScratchMemory_l160_115;
  wire                when_BankedScratchMemory_l160_116;
  wire                when_BankedScratchMemory_l160_117;
  wire                when_BankedScratchMemory_l160_118;
  wire                when_BankedScratchMemory_l160_119;
  wire       [2:0]    _zz_when_BankedScratchMemory_l160_15;
  wire       [7:0]    _zz_io_reads_1_addr_7;
  reg        [31:0]   _zz_io_valuReadData_1_7;
  wire                when_BankedScratchMemory_l160_120;
  wire                when_BankedScratchMemory_l160_121;
  wire                when_BankedScratchMemory_l160_122;
  wire                when_BankedScratchMemory_l160_123;
  wire                when_BankedScratchMemory_l160_124;
  wire                when_BankedScratchMemory_l160_125;
  wire                when_BankedScratchMemory_l160_126;
  wire                when_BankedScratchMemory_l160_127;
  wire       [2:0]    scalarBankReq_0;
  wire       [2:0]    scalarBankReq_1;
  wire       [2:0]    scalarBankReq_2;
  wire       [2:0]    scalarBankReq_3;
  wire       [2:0]    scalarBankReq_4;
  wire       [2:0]    scalarBankReq_5;
  wire       [2:0]    scalarBankReq_6;
  wire       [2:0]    scalarBankReq_7;
  wire       [2:0]    scalarBankReq_8;
  wire       [7:0]    scalarBankRow_0;
  wire       [7:0]    scalarBankRow_1;
  wire       [7:0]    scalarBankRow_2;
  wire       [7:0]    scalarBankRow_3;
  wire       [7:0]    scalarBankRow_4;
  wire       [7:0]    scalarBankRow_5;
  wire       [7:0]    scalarBankRow_6;
  wire       [7:0]    scalarBankRow_7;
  wire       [7:0]    scalarBankRow_8;
  wire                _zz_when_BankedScratchMemory_l203;
  wire                when_BankedScratchMemory_l203;
  wire                when_BankedScratchMemory_l206;
  wire                when_BankedScratchMemory_l206_1;
  wire                when_BankedScratchMemory_l206_2;
  wire                when_BankedScratchMemory_l206_3;
  wire                when_BankedScratchMemory_l206_4;
  wire                when_BankedScratchMemory_l206_5;
  wire                when_BankedScratchMemory_l206_6;
  wire                when_BankedScratchMemory_l206_7;
  wire                when_BankedScratchMemory_l213;
  wire                _zz_when_BankedScratchMemory_l203_1;
  wire                when_BankedScratchMemory_l203_1;
  wire                when_BankedScratchMemory_l206_8;
  wire                when_BankedScratchMemory_l206_9;
  wire                when_BankedScratchMemory_l206_10;
  wire                when_BankedScratchMemory_l206_11;
  wire                when_BankedScratchMemory_l206_12;
  wire                when_BankedScratchMemory_l206_13;
  wire                when_BankedScratchMemory_l206_14;
  wire                when_BankedScratchMemory_l206_15;
  wire                when_BankedScratchMemory_l213_1;
  wire                _zz_when_BankedScratchMemory_l203_2;
  wire                when_BankedScratchMemory_l203_2;
  wire                when_BankedScratchMemory_l206_16;
  wire                when_BankedScratchMemory_l206_17;
  wire                when_BankedScratchMemory_l206_18;
  wire                when_BankedScratchMemory_l206_19;
  wire                when_BankedScratchMemory_l206_20;
  wire                when_BankedScratchMemory_l206_21;
  wire                when_BankedScratchMemory_l206_22;
  wire                when_BankedScratchMemory_l206_23;
  wire                when_BankedScratchMemory_l213_2;
  wire                _zz_when_BankedScratchMemory_l203_3;
  wire                when_BankedScratchMemory_l203_3;
  wire                when_BankedScratchMemory_l206_24;
  wire                when_BankedScratchMemory_l206_25;
  wire                when_BankedScratchMemory_l206_26;
  wire                when_BankedScratchMemory_l206_27;
  wire                when_BankedScratchMemory_l206_28;
  wire                when_BankedScratchMemory_l206_29;
  wire                when_BankedScratchMemory_l206_30;
  wire                when_BankedScratchMemory_l206_31;
  wire                when_BankedScratchMemory_l213_3;
  wire                _zz_when_BankedScratchMemory_l203_4;
  wire                when_BankedScratchMemory_l203_4;
  wire                when_BankedScratchMemory_l206_32;
  wire                when_BankedScratchMemory_l206_33;
  wire                when_BankedScratchMemory_l206_34;
  wire                when_BankedScratchMemory_l206_35;
  wire                when_BankedScratchMemory_l206_36;
  wire                when_BankedScratchMemory_l206_37;
  wire                when_BankedScratchMemory_l206_38;
  wire                when_BankedScratchMemory_l206_39;
  wire                when_BankedScratchMemory_l213_4;
  wire                _zz_when_BankedScratchMemory_l203_5;
  wire                when_BankedScratchMemory_l203_5;
  wire                when_BankedScratchMemory_l206_40;
  wire                when_BankedScratchMemory_l206_41;
  wire                when_BankedScratchMemory_l206_42;
  wire                when_BankedScratchMemory_l206_43;
  wire                when_BankedScratchMemory_l206_44;
  wire                when_BankedScratchMemory_l206_45;
  wire                when_BankedScratchMemory_l206_46;
  wire                when_BankedScratchMemory_l206_47;
  wire                when_BankedScratchMemory_l213_5;
  wire                _zz_when_BankedScratchMemory_l203_6;
  wire                when_BankedScratchMemory_l203_6;
  wire                when_BankedScratchMemory_l206_48;
  wire                when_BankedScratchMemory_l206_49;
  wire                when_BankedScratchMemory_l206_50;
  wire                when_BankedScratchMemory_l206_51;
  wire                when_BankedScratchMemory_l206_52;
  wire                when_BankedScratchMemory_l206_53;
  wire                when_BankedScratchMemory_l206_54;
  wire                when_BankedScratchMemory_l206_55;
  wire                when_BankedScratchMemory_l213_6;
  wire                _zz_when_BankedScratchMemory_l203_7;
  wire                when_BankedScratchMemory_l203_7;
  wire                when_BankedScratchMemory_l206_56;
  wire                when_BankedScratchMemory_l206_57;
  wire                when_BankedScratchMemory_l206_58;
  wire                when_BankedScratchMemory_l206_59;
  wire                when_BankedScratchMemory_l206_60;
  wire                when_BankedScratchMemory_l206_61;
  wire                when_BankedScratchMemory_l206_62;
  wire                when_BankedScratchMemory_l206_63;
  wire                when_BankedScratchMemory_l213_7;
  wire                _zz_when_BankedScratchMemory_l203_8;
  wire                when_BankedScratchMemory_l203_8;
  wire                when_BankedScratchMemory_l206_64;
  wire                when_BankedScratchMemory_l206_65;
  wire                when_BankedScratchMemory_l206_66;
  wire                when_BankedScratchMemory_l206_67;
  wire                when_BankedScratchMemory_l206_68;
  wire                when_BankedScratchMemory_l206_69;
  wire                when_BankedScratchMemory_l206_70;
  wire                when_BankedScratchMemory_l206_71;
  wire                when_BankedScratchMemory_l213_8;
  wire                when_BankedScratchMemory_l222;
  wire                when_BankedScratchMemory_l222_1;
  wire                when_BankedScratchMemory_l222_2;
  wire                when_BankedScratchMemory_l222_3;
  wire                when_BankedScratchMemory_l222_4;
  wire                when_BankedScratchMemory_l222_5;
  wire                when_BankedScratchMemory_l222_6;
  wire                when_BankedScratchMemory_l222_7;
  wire                when_BankedScratchMemory_l222_8;
  wire                when_BankedScratchMemory_l222_9;
  wire                when_BankedScratchMemory_l222_10;
  wire                when_BankedScratchMemory_l222_11;
  wire                when_BankedScratchMemory_l222_12;
  wire                when_BankedScratchMemory_l222_13;
  wire                when_BankedScratchMemory_l222_14;
  wire                when_BankedScratchMemory_l222_15;
  wire                when_BankedScratchMemory_l222_16;
  wire                when_BankedScratchMemory_l222_17;
  wire                when_BankedScratchMemory_l222_18;
  wire                when_BankedScratchMemory_l222_19;
  wire                when_BankedScratchMemory_l222_20;
  wire                when_BankedScratchMemory_l222_21;
  wire                when_BankedScratchMemory_l222_22;
  wire                when_BankedScratchMemory_l222_23;
  wire                when_BankedScratchMemory_l222_24;
  wire                when_BankedScratchMemory_l222_25;
  wire                when_BankedScratchMemory_l222_26;
  wire                when_BankedScratchMemory_l222_27;
  wire                when_BankedScratchMemory_l222_28;
  wire                when_BankedScratchMemory_l222_29;
  wire                when_BankedScratchMemory_l222_30;
  wire                when_BankedScratchMemory_l222_31;
  wire                when_BankedScratchMemory_l222_32;
  wire                when_BankedScratchMemory_l222_33;
  wire                when_BankedScratchMemory_l222_34;
  wire                when_BankedScratchMemory_l222_35;
  wire                when_BankedScratchMemory_l222_36;
  wire                when_BankedScratchMemory_l222_37;
  wire                when_BankedScratchMemory_l222_38;
  wire                when_BankedScratchMemory_l222_39;
  wire                when_BankedScratchMemory_l222_40;
  wire                when_BankedScratchMemory_l222_41;
  wire                when_BankedScratchMemory_l222_42;
  wire                when_BankedScratchMemory_l222_43;
  wire                when_BankedScratchMemory_l222_44;
  wire                when_BankedScratchMemory_l222_45;
  wire                when_BankedScratchMemory_l222_46;
  wire                when_BankedScratchMemory_l222_47;
  wire                when_BankedScratchMemory_l222_48;
  wire                when_BankedScratchMemory_l222_49;
  wire                when_BankedScratchMemory_l222_50;
  wire                when_BankedScratchMemory_l222_51;
  wire                when_BankedScratchMemory_l222_52;
  wire                when_BankedScratchMemory_l222_53;
  wire                when_BankedScratchMemory_l222_54;
  wire                when_BankedScratchMemory_l222_55;
  wire                when_BankedScratchMemory_l222_56;
  wire                when_BankedScratchMemory_l222_57;
  wire                when_BankedScratchMemory_l222_58;
  wire                when_BankedScratchMemory_l222_59;
  wire                when_BankedScratchMemory_l222_60;
  wire                when_BankedScratchMemory_l222_61;
  wire                when_BankedScratchMemory_l222_62;
  wire                when_BankedScratchMemory_l222_63;
  wire                when_BankedScratchMemory_l222_64;
  wire                when_BankedScratchMemory_l222_65;
  wire                when_BankedScratchMemory_l222_66;
  wire                when_BankedScratchMemory_l222_67;
  wire                when_BankedScratchMemory_l222_68;
  wire                when_BankedScratchMemory_l222_69;
  wire                when_BankedScratchMemory_l222_70;
  wire                when_BankedScratchMemory_l222_71;
  wire       [2:0]    _zz_when_BankedScratchMemory_l242;
  wire       [7:0]    _zz_io_write_addr;
  wire                when_BankedScratchMemory_l242;
  wire                when_BankedScratchMemory_l242_1;
  wire                when_BankedScratchMemory_l242_2;
  wire                when_BankedScratchMemory_l242_3;
  wire                when_BankedScratchMemory_l242_4;
  wire                when_BankedScratchMemory_l242_5;
  wire                when_BankedScratchMemory_l242_6;
  wire                when_BankedScratchMemory_l242_7;
  wire       [2:0]    _zz_when_BankedScratchMemory_l242_1;
  wire       [7:0]    _zz_io_write_addr_1;
  wire                when_BankedScratchMemory_l242_8;
  wire                when_BankedScratchMemory_l242_9;
  wire                when_BankedScratchMemory_l242_10;
  wire                when_BankedScratchMemory_l242_11;
  wire                when_BankedScratchMemory_l242_12;
  wire                when_BankedScratchMemory_l242_13;
  wire                when_BankedScratchMemory_l242_14;
  wire                when_BankedScratchMemory_l242_15;
  wire       [2:0]    _zz_when_BankedScratchMemory_l242_2;
  wire       [7:0]    _zz_io_write_addr_2;
  wire                when_BankedScratchMemory_l242_16;
  wire                when_BankedScratchMemory_l242_17;
  wire                when_BankedScratchMemory_l242_18;
  wire                when_BankedScratchMemory_l242_19;
  wire                when_BankedScratchMemory_l242_20;
  wire                when_BankedScratchMemory_l242_21;
  wire                when_BankedScratchMemory_l242_22;
  wire                when_BankedScratchMemory_l242_23;
  wire       [2:0]    _zz_when_BankedScratchMemory_l242_3;
  wire       [7:0]    _zz_io_write_addr_3;
  wire                when_BankedScratchMemory_l242_24;
  wire                when_BankedScratchMemory_l242_25;
  wire                when_BankedScratchMemory_l242_26;
  wire                when_BankedScratchMemory_l242_27;
  wire                when_BankedScratchMemory_l242_28;
  wire                when_BankedScratchMemory_l242_29;
  wire                when_BankedScratchMemory_l242_30;
  wire                when_BankedScratchMemory_l242_31;
  wire       [2:0]    _zz_when_BankedScratchMemory_l242_4;
  wire       [7:0]    _zz_io_write_addr_4;
  wire                when_BankedScratchMemory_l242_32;
  wire                when_BankedScratchMemory_l242_33;
  wire                when_BankedScratchMemory_l242_34;
  wire                when_BankedScratchMemory_l242_35;
  wire                when_BankedScratchMemory_l242_36;
  wire                when_BankedScratchMemory_l242_37;
  wire                when_BankedScratchMemory_l242_38;
  wire                when_BankedScratchMemory_l242_39;
  wire       [2:0]    _zz_when_BankedScratchMemory_l242_5;
  wire       [7:0]    _zz_io_write_addr_5;
  wire                when_BankedScratchMemory_l242_40;
  wire                when_BankedScratchMemory_l242_41;
  wire                when_BankedScratchMemory_l242_42;
  wire                when_BankedScratchMemory_l242_43;
  wire                when_BankedScratchMemory_l242_44;
  wire                when_BankedScratchMemory_l242_45;
  wire                when_BankedScratchMemory_l242_46;
  wire                when_BankedScratchMemory_l242_47;
  wire       [2:0]    _zz_when_BankedScratchMemory_l242_6;
  wire       [7:0]    _zz_io_write_addr_6;
  wire                when_BankedScratchMemory_l242_48;
  wire                when_BankedScratchMemory_l242_49;
  wire                when_BankedScratchMemory_l242_50;
  wire                when_BankedScratchMemory_l242_51;
  wire                when_BankedScratchMemory_l242_52;
  wire                when_BankedScratchMemory_l242_53;
  wire                when_BankedScratchMemory_l242_54;
  wire                when_BankedScratchMemory_l242_55;
  wire       [2:0]    _zz_when_BankedScratchMemory_l242_7;
  wire       [7:0]    _zz_io_write_addr_7;
  wire                when_BankedScratchMemory_l242_56;
  wire                when_BankedScratchMemory_l242_57;
  wire                when_BankedScratchMemory_l242_58;
  wire                when_BankedScratchMemory_l242_59;
  wire                when_BankedScratchMemory_l242_60;
  wire                when_BankedScratchMemory_l242_61;
  wire                when_BankedScratchMemory_l242_62;
  wire                when_BankedScratchMemory_l242_63;
  wire       [2:0]    _zz_when_BankedScratchMemory_l242_8;
  wire       [7:0]    _zz_io_write_addr_8;
  wire                when_BankedScratchMemory_l242_64;
  wire                when_BankedScratchMemory_l242_65;
  wire                when_BankedScratchMemory_l242_66;
  wire                when_BankedScratchMemory_l242_67;
  wire                when_BankedScratchMemory_l242_68;
  wire                when_BankedScratchMemory_l242_69;
  wire                when_BankedScratchMemory_l242_70;
  wire                when_BankedScratchMemory_l242_71;
  wire       [2:0]    _zz_when_BankedScratchMemory_l242_9;
  wire       [7:0]    _zz_io_write_addr_9;
  wire                when_BankedScratchMemory_l242_72;
  wire                when_BankedScratchMemory_l242_73;
  wire                when_BankedScratchMemory_l242_74;
  wire                when_BankedScratchMemory_l242_75;
  wire                when_BankedScratchMemory_l242_76;
  wire                when_BankedScratchMemory_l242_77;
  wire                when_BankedScratchMemory_l242_78;
  wire                when_BankedScratchMemory_l242_79;
  wire       [2:0]    _zz_when_BankedScratchMemory_l242_10;
  wire       [7:0]    _zz_io_write_addr_10;
  wire                when_BankedScratchMemory_l242_80;
  wire                when_BankedScratchMemory_l242_81;
  wire                when_BankedScratchMemory_l242_82;
  wire                when_BankedScratchMemory_l242_83;
  wire                when_BankedScratchMemory_l242_84;
  wire                when_BankedScratchMemory_l242_85;
  wire                when_BankedScratchMemory_l242_86;
  wire                when_BankedScratchMemory_l242_87;
  wire       [2:0]    _zz_when_BankedScratchMemory_l242_11;
  wire       [7:0]    _zz_io_write_addr_11;
  wire                when_BankedScratchMemory_l242_88;
  wire                when_BankedScratchMemory_l242_89;
  wire                when_BankedScratchMemory_l242_90;
  wire                when_BankedScratchMemory_l242_91;
  wire                when_BankedScratchMemory_l242_92;
  wire                when_BankedScratchMemory_l242_93;
  wire                when_BankedScratchMemory_l242_94;
  wire                when_BankedScratchMemory_l242_95;
  wire       [2:0]    _zz_when_BankedScratchMemory_l242_12;
  wire       [7:0]    _zz_io_write_addr_12;
  wire                when_BankedScratchMemory_l242_96;
  wire                when_BankedScratchMemory_l242_97;
  wire                when_BankedScratchMemory_l242_98;
  wire                when_BankedScratchMemory_l242_99;
  wire                when_BankedScratchMemory_l242_100;
  wire                when_BankedScratchMemory_l242_101;
  wire                when_BankedScratchMemory_l242_102;
  wire                when_BankedScratchMemory_l242_103;
  wire       [2:0]    _zz_when_BankedScratchMemory_l242_13;
  wire       [7:0]    _zz_io_write_addr_13;
  wire                when_BankedScratchMemory_l242_104;
  wire                when_BankedScratchMemory_l242_105;
  wire                when_BankedScratchMemory_l242_106;
  wire                when_BankedScratchMemory_l242_107;
  wire                when_BankedScratchMemory_l242_108;
  wire                when_BankedScratchMemory_l242_109;
  wire                when_BankedScratchMemory_l242_110;
  wire                when_BankedScratchMemory_l242_111;
  wire       [2:0]    _zz_when_BankedScratchMemory_l242_14;
  wire       [7:0]    _zz_io_write_addr_14;
  wire                when_BankedScratchMemory_l242_112;
  wire                when_BankedScratchMemory_l242_113;
  wire                when_BankedScratchMemory_l242_114;
  wire                when_BankedScratchMemory_l242_115;
  wire                when_BankedScratchMemory_l242_116;
  wire                when_BankedScratchMemory_l242_117;
  wire                when_BankedScratchMemory_l242_118;
  wire                when_BankedScratchMemory_l242_119;
  wire       [2:0]    _zz_when_BankedScratchMemory_l242_15;
  wire       [7:0]    _zz_io_write_addr_15;
  wire                when_BankedScratchMemory_l242_120;
  wire                when_BankedScratchMemory_l242_121;
  wire                when_BankedScratchMemory_l242_122;
  wire                when_BankedScratchMemory_l242_123;
  wire                when_BankedScratchMemory_l242_124;
  wire                when_BankedScratchMemory_l242_125;
  wire                when_BankedScratchMemory_l242_126;
  wire                when_BankedScratchMemory_l242_127;
  wire       [2:0]    _zz_when_BankedScratchMemory_l242_16;
  wire       [7:0]    _zz_io_write_addr_16;
  wire                when_BankedScratchMemory_l242_128;
  wire                when_BankedScratchMemory_l242_129;
  wire                when_BankedScratchMemory_l242_130;
  wire                when_BankedScratchMemory_l242_131;
  wire                when_BankedScratchMemory_l242_132;
  wire                when_BankedScratchMemory_l242_133;
  wire                when_BankedScratchMemory_l242_134;
  wire                when_BankedScratchMemory_l242_135;
  wire       [2:0]    _zz_when_BankedScratchMemory_l242_17;
  wire       [7:0]    _zz_io_write_addr_17;
  wire                when_BankedScratchMemory_l242_136;
  wire                when_BankedScratchMemory_l242_137;
  wire                when_BankedScratchMemory_l242_138;
  wire                when_BankedScratchMemory_l242_139;
  wire                when_BankedScratchMemory_l242_140;
  wire                when_BankedScratchMemory_l242_141;
  wire                when_BankedScratchMemory_l242_142;
  wire                when_BankedScratchMemory_l242_143;
  wire       [2:0]    _zz_when_BankedScratchMemory_l242_18;
  wire       [7:0]    _zz_io_write_addr_18;
  wire                when_BankedScratchMemory_l242_144;
  wire                when_BankedScratchMemory_l242_145;
  wire                when_BankedScratchMemory_l242_146;
  wire                when_BankedScratchMemory_l242_147;
  wire                when_BankedScratchMemory_l242_148;
  wire                when_BankedScratchMemory_l242_149;
  wire                when_BankedScratchMemory_l242_150;
  wire                when_BankedScratchMemory_l242_151;
  wire       [2:0]    _zz_when_BankedScratchMemory_l242_19;
  wire       [7:0]    _zz_io_write_addr_19;
  wire                when_BankedScratchMemory_l242_152;
  wire                when_BankedScratchMemory_l242_153;
  wire                when_BankedScratchMemory_l242_154;
  wire                when_BankedScratchMemory_l242_155;
  wire                when_BankedScratchMemory_l242_156;
  wire                when_BankedScratchMemory_l242_157;
  wire                when_BankedScratchMemory_l242_158;
  wire                when_BankedScratchMemory_l242_159;
  wire       [2:0]    _zz_when_BankedScratchMemory_l242_20;
  wire       [7:0]    _zz_io_write_addr_20;
  wire                when_BankedScratchMemory_l242_160;
  wire                when_BankedScratchMemory_l242_161;
  wire                when_BankedScratchMemory_l242_162;
  wire                when_BankedScratchMemory_l242_163;
  wire                when_BankedScratchMemory_l242_164;
  wire                when_BankedScratchMemory_l242_165;
  wire                when_BankedScratchMemory_l242_166;
  wire                when_BankedScratchMemory_l242_167;
  wire       [2:0]    _zz_when_BankedScratchMemory_l242_21;
  wire       [7:0]    _zz_io_write_addr_21;
  wire                when_BankedScratchMemory_l242_168;
  wire                when_BankedScratchMemory_l242_169;
  wire                when_BankedScratchMemory_l242_170;
  wire                when_BankedScratchMemory_l242_171;
  wire                when_BankedScratchMemory_l242_172;
  wire                when_BankedScratchMemory_l242_173;
  wire                when_BankedScratchMemory_l242_174;
  wire                when_BankedScratchMemory_l242_175;
  wire       [2:0]    _zz_when_BankedScratchMemory_l242_22;
  wire       [7:0]    _zz_io_write_addr_22;
  wire                when_BankedScratchMemory_l242_176;
  wire                when_BankedScratchMemory_l242_177;
  wire                when_BankedScratchMemory_l242_178;
  wire                when_BankedScratchMemory_l242_179;
  wire                when_BankedScratchMemory_l242_180;
  wire                when_BankedScratchMemory_l242_181;
  wire                when_BankedScratchMemory_l242_182;
  wire                when_BankedScratchMemory_l242_183;
  wire       [2:0]    _zz_when_BankedScratchMemory_l242_23;
  wire       [7:0]    _zz_io_write_addr_23;
  wire                when_BankedScratchMemory_l242_184;
  wire                when_BankedScratchMemory_l242_185;
  wire                when_BankedScratchMemory_l242_186;
  wire                when_BankedScratchMemory_l242_187;
  wire                when_BankedScratchMemory_l242_188;
  wire                when_BankedScratchMemory_l242_189;
  wire                when_BankedScratchMemory_l242_190;
  wire                when_BankedScratchMemory_l242_191;
  wire       [2:0]    _zz_when_BankedScratchMemory_l242_24;
  wire       [7:0]    _zz_io_write_addr_24;
  wire                when_BankedScratchMemory_l242_192;
  wire                when_BankedScratchMemory_l242_193;
  wire                when_BankedScratchMemory_l242_194;
  wire                when_BankedScratchMemory_l242_195;
  wire                when_BankedScratchMemory_l242_196;
  wire                when_BankedScratchMemory_l242_197;
  wire                when_BankedScratchMemory_l242_198;
  wire                when_BankedScratchMemory_l242_199;
  wire       [2:0]    _zz_when_BankedScratchMemory_l242_25;
  wire       [7:0]    _zz_io_write_addr_25;
  wire                when_BankedScratchMemory_l242_200;
  wire                when_BankedScratchMemory_l242_201;
  wire                when_BankedScratchMemory_l242_202;
  wire                when_BankedScratchMemory_l242_203;
  wire                when_BankedScratchMemory_l242_204;
  wire                when_BankedScratchMemory_l242_205;
  wire                when_BankedScratchMemory_l242_206;
  wire                when_BankedScratchMemory_l242_207;
  wire       [2:0]    _zz_when_BankedScratchMemory_l242_26;
  wire       [7:0]    _zz_io_write_addr_26;
  wire                when_BankedScratchMemory_l242_208;
  wire                when_BankedScratchMemory_l242_209;
  wire                when_BankedScratchMemory_l242_210;
  wire                when_BankedScratchMemory_l242_211;
  wire                when_BankedScratchMemory_l242_212;
  wire                when_BankedScratchMemory_l242_213;
  wire                when_BankedScratchMemory_l242_214;
  wire                when_BankedScratchMemory_l242_215;
  wire       [2:0]    _zz_when_BankedScratchMemory_l242_27;
  wire       [7:0]    _zz_io_write_addr_27;
  wire                when_BankedScratchMemory_l242_216;
  wire                when_BankedScratchMemory_l242_217;
  wire                when_BankedScratchMemory_l242_218;
  wire                when_BankedScratchMemory_l242_219;
  wire                when_BankedScratchMemory_l242_220;
  wire                when_BankedScratchMemory_l242_221;
  wire                when_BankedScratchMemory_l242_222;
  wire                when_BankedScratchMemory_l242_223;

  assign _zz__zz_when_BankedScratchMemory_l203_7 = (scalarBankReq_0 == scalarBankReq_7);
  assign _zz__zz_when_BankedScratchMemory_l203_7_1 = (scalarBankReq_1 == scalarBankReq_7);
  assign _zz__zz_when_BankedScratchMemory_l203_8 = (io_scalarReadEn_0 && (scalarBankReq_0 == scalarBankReq_8));
  assign _zz__zz_when_BankedScratchMemory_l203_8_1 = (io_scalarReadEn_1 && (scalarBankReq_1 == scalarBankReq_8));
  assign _zz__zz_when_BankedScratchMemory_l203_8_2 = (scalarBankReq_2 == scalarBankReq_8);
  ScratchBank banks_0 (
    .io_reads_0_addr (banks_0_io_reads_0_addr[7:0] ), //i
    .io_reads_0_en   (banks_0_io_reads_0_en        ), //i
    .io_reads_0_data (banks_0_io_reads_0_data[31:0]), //o
    .io_reads_1_addr (banks_0_io_reads_1_addr[7:0] ), //i
    .io_reads_1_en   (banks_0_io_reads_1_en        ), //i
    .io_reads_1_data (banks_0_io_reads_1_data[31:0]), //o
    .io_reads_2_addr (banks_0_io_reads_2_addr[7:0] ), //i
    .io_reads_2_en   (banks_0_io_reads_2_en        ), //i
    .io_reads_2_data (banks_0_io_reads_2_data[31:0]), //o
    .io_write_addr   (banks_0_io_write_addr[7:0]   ), //i
    .io_write_data   (banks_0_io_write_data[31:0]  ), //i
    .io_write_en     (banks_0_io_write_en          ), //i
    .clk             (clk                          ), //i
    .reset           (reset                        )  //i
  );
  ScratchBank banks_1 (
    .io_reads_0_addr (banks_1_io_reads_0_addr[7:0] ), //i
    .io_reads_0_en   (banks_1_io_reads_0_en        ), //i
    .io_reads_0_data (banks_1_io_reads_0_data[31:0]), //o
    .io_reads_1_addr (banks_1_io_reads_1_addr[7:0] ), //i
    .io_reads_1_en   (banks_1_io_reads_1_en        ), //i
    .io_reads_1_data (banks_1_io_reads_1_data[31:0]), //o
    .io_reads_2_addr (banks_1_io_reads_2_addr[7:0] ), //i
    .io_reads_2_en   (banks_1_io_reads_2_en        ), //i
    .io_reads_2_data (banks_1_io_reads_2_data[31:0]), //o
    .io_write_addr   (banks_1_io_write_addr[7:0]   ), //i
    .io_write_data   (banks_1_io_write_data[31:0]  ), //i
    .io_write_en     (banks_1_io_write_en          ), //i
    .clk             (clk                          ), //i
    .reset           (reset                        )  //i
  );
  ScratchBank banks_2 (
    .io_reads_0_addr (banks_2_io_reads_0_addr[7:0] ), //i
    .io_reads_0_en   (banks_2_io_reads_0_en        ), //i
    .io_reads_0_data (banks_2_io_reads_0_data[31:0]), //o
    .io_reads_1_addr (banks_2_io_reads_1_addr[7:0] ), //i
    .io_reads_1_en   (banks_2_io_reads_1_en        ), //i
    .io_reads_1_data (banks_2_io_reads_1_data[31:0]), //o
    .io_reads_2_addr (banks_2_io_reads_2_addr[7:0] ), //i
    .io_reads_2_en   (banks_2_io_reads_2_en        ), //i
    .io_reads_2_data (banks_2_io_reads_2_data[31:0]), //o
    .io_write_addr   (banks_2_io_write_addr[7:0]   ), //i
    .io_write_data   (banks_2_io_write_data[31:0]  ), //i
    .io_write_en     (banks_2_io_write_en          ), //i
    .clk             (clk                          ), //i
    .reset           (reset                        )  //i
  );
  ScratchBank banks_3 (
    .io_reads_0_addr (banks_3_io_reads_0_addr[7:0] ), //i
    .io_reads_0_en   (banks_3_io_reads_0_en        ), //i
    .io_reads_0_data (banks_3_io_reads_0_data[31:0]), //o
    .io_reads_1_addr (banks_3_io_reads_1_addr[7:0] ), //i
    .io_reads_1_en   (banks_3_io_reads_1_en        ), //i
    .io_reads_1_data (banks_3_io_reads_1_data[31:0]), //o
    .io_reads_2_addr (banks_3_io_reads_2_addr[7:0] ), //i
    .io_reads_2_en   (banks_3_io_reads_2_en        ), //i
    .io_reads_2_data (banks_3_io_reads_2_data[31:0]), //o
    .io_write_addr   (banks_3_io_write_addr[7:0]   ), //i
    .io_write_data   (banks_3_io_write_data[31:0]  ), //i
    .io_write_en     (banks_3_io_write_en          ), //i
    .clk             (clk                          ), //i
    .reset           (reset                        )  //i
  );
  ScratchBank banks_4 (
    .io_reads_0_addr (banks_4_io_reads_0_addr[7:0] ), //i
    .io_reads_0_en   (banks_4_io_reads_0_en        ), //i
    .io_reads_0_data (banks_4_io_reads_0_data[31:0]), //o
    .io_reads_1_addr (banks_4_io_reads_1_addr[7:0] ), //i
    .io_reads_1_en   (banks_4_io_reads_1_en        ), //i
    .io_reads_1_data (banks_4_io_reads_1_data[31:0]), //o
    .io_reads_2_addr (banks_4_io_reads_2_addr[7:0] ), //i
    .io_reads_2_en   (banks_4_io_reads_2_en        ), //i
    .io_reads_2_data (banks_4_io_reads_2_data[31:0]), //o
    .io_write_addr   (banks_4_io_write_addr[7:0]   ), //i
    .io_write_data   (banks_4_io_write_data[31:0]  ), //i
    .io_write_en     (banks_4_io_write_en          ), //i
    .clk             (clk                          ), //i
    .reset           (reset                        )  //i
  );
  ScratchBank banks_5 (
    .io_reads_0_addr (banks_5_io_reads_0_addr[7:0] ), //i
    .io_reads_0_en   (banks_5_io_reads_0_en        ), //i
    .io_reads_0_data (banks_5_io_reads_0_data[31:0]), //o
    .io_reads_1_addr (banks_5_io_reads_1_addr[7:0] ), //i
    .io_reads_1_en   (banks_5_io_reads_1_en        ), //i
    .io_reads_1_data (banks_5_io_reads_1_data[31:0]), //o
    .io_reads_2_addr (banks_5_io_reads_2_addr[7:0] ), //i
    .io_reads_2_en   (banks_5_io_reads_2_en        ), //i
    .io_reads_2_data (banks_5_io_reads_2_data[31:0]), //o
    .io_write_addr   (banks_5_io_write_addr[7:0]   ), //i
    .io_write_data   (banks_5_io_write_data[31:0]  ), //i
    .io_write_en     (banks_5_io_write_en          ), //i
    .clk             (clk                          ), //i
    .reset           (reset                        )  //i
  );
  ScratchBank banks_6 (
    .io_reads_0_addr (banks_6_io_reads_0_addr[7:0] ), //i
    .io_reads_0_en   (banks_6_io_reads_0_en        ), //i
    .io_reads_0_data (banks_6_io_reads_0_data[31:0]), //o
    .io_reads_1_addr (banks_6_io_reads_1_addr[7:0] ), //i
    .io_reads_1_en   (banks_6_io_reads_1_en        ), //i
    .io_reads_1_data (banks_6_io_reads_1_data[31:0]), //o
    .io_reads_2_addr (banks_6_io_reads_2_addr[7:0] ), //i
    .io_reads_2_en   (banks_6_io_reads_2_en        ), //i
    .io_reads_2_data (banks_6_io_reads_2_data[31:0]), //o
    .io_write_addr   (banks_6_io_write_addr[7:0]   ), //i
    .io_write_data   (banks_6_io_write_data[31:0]  ), //i
    .io_write_en     (banks_6_io_write_en          ), //i
    .clk             (clk                          ), //i
    .reset           (reset                        )  //i
  );
  ScratchBank banks_7 (
    .io_reads_0_addr (banks_7_io_reads_0_addr[7:0] ), //i
    .io_reads_0_en   (banks_7_io_reads_0_en        ), //i
    .io_reads_0_data (banks_7_io_reads_0_data[31:0]), //o
    .io_reads_1_addr (banks_7_io_reads_1_addr[7:0] ), //i
    .io_reads_1_en   (banks_7_io_reads_1_en        ), //i
    .io_reads_1_data (banks_7_io_reads_1_data[31:0]), //o
    .io_reads_2_addr (banks_7_io_reads_2_addr[7:0] ), //i
    .io_reads_2_en   (banks_7_io_reads_2_en        ), //i
    .io_reads_2_data (banks_7_io_reads_2_data[31:0]), //o
    .io_write_addr   (banks_7_io_write_addr[7:0]   ), //i
    .io_write_data   (banks_7_io_write_data[31:0]  ), //i
    .io_write_en     (banks_7_io_write_en          ), //i
    .clk             (clk                          ), //i
    .reset           (reset                        )  //i
  );
  always @(*) begin
    banks_0_io_reads_0_addr = 8'h0;
    if(when_BankedScratchMemory_l160) begin
      banks_0_io_reads_0_addr = _zz_io_reads_0_addr;
    end
    if(when_BankedScratchMemory_l160_8) begin
      banks_0_io_reads_0_addr = _zz_io_reads_0_addr_1;
    end
    if(when_BankedScratchMemory_l160_16) begin
      banks_0_io_reads_0_addr = _zz_io_reads_0_addr_2;
    end
    if(when_BankedScratchMemory_l160_24) begin
      banks_0_io_reads_0_addr = _zz_io_reads_0_addr_3;
    end
    if(when_BankedScratchMemory_l160_32) begin
      banks_0_io_reads_0_addr = _zz_io_reads_0_addr_4;
    end
    if(when_BankedScratchMemory_l160_40) begin
      banks_0_io_reads_0_addr = _zz_io_reads_0_addr_5;
    end
    if(when_BankedScratchMemory_l160_48) begin
      banks_0_io_reads_0_addr = _zz_io_reads_0_addr_6;
    end
    if(when_BankedScratchMemory_l160_56) begin
      banks_0_io_reads_0_addr = _zz_io_reads_0_addr_7;
    end
  end

  always @(*) begin
    banks_0_io_reads_0_en = 1'b0;
    if(when_BankedScratchMemory_l160) begin
      banks_0_io_reads_0_en = io_valuReadEn_0_0;
    end
    if(when_BankedScratchMemory_l160_8) begin
      banks_0_io_reads_0_en = io_valuReadEn_0_1;
    end
    if(when_BankedScratchMemory_l160_16) begin
      banks_0_io_reads_0_en = io_valuReadEn_0_2;
    end
    if(when_BankedScratchMemory_l160_24) begin
      banks_0_io_reads_0_en = io_valuReadEn_0_3;
    end
    if(when_BankedScratchMemory_l160_32) begin
      banks_0_io_reads_0_en = io_valuReadEn_0_4;
    end
    if(when_BankedScratchMemory_l160_40) begin
      banks_0_io_reads_0_en = io_valuReadEn_0_5;
    end
    if(when_BankedScratchMemory_l160_48) begin
      banks_0_io_reads_0_en = io_valuReadEn_0_6;
    end
    if(when_BankedScratchMemory_l160_56) begin
      banks_0_io_reads_0_en = io_valuReadEn_0_7;
    end
  end

  always @(*) begin
    banks_0_io_reads_1_addr = 8'h0;
    if(when_BankedScratchMemory_l160_64) begin
      banks_0_io_reads_1_addr = _zz_io_reads_1_addr;
    end
    if(when_BankedScratchMemory_l160_72) begin
      banks_0_io_reads_1_addr = _zz_io_reads_1_addr_1;
    end
    if(when_BankedScratchMemory_l160_80) begin
      banks_0_io_reads_1_addr = _zz_io_reads_1_addr_2;
    end
    if(when_BankedScratchMemory_l160_88) begin
      banks_0_io_reads_1_addr = _zz_io_reads_1_addr_3;
    end
    if(when_BankedScratchMemory_l160_96) begin
      banks_0_io_reads_1_addr = _zz_io_reads_1_addr_4;
    end
    if(when_BankedScratchMemory_l160_104) begin
      banks_0_io_reads_1_addr = _zz_io_reads_1_addr_5;
    end
    if(when_BankedScratchMemory_l160_112) begin
      banks_0_io_reads_1_addr = _zz_io_reads_1_addr_6;
    end
    if(when_BankedScratchMemory_l160_120) begin
      banks_0_io_reads_1_addr = _zz_io_reads_1_addr_7;
    end
  end

  always @(*) begin
    banks_0_io_reads_1_en = 1'b0;
    if(when_BankedScratchMemory_l160_64) begin
      banks_0_io_reads_1_en = io_valuReadEn_1_0;
    end
    if(when_BankedScratchMemory_l160_72) begin
      banks_0_io_reads_1_en = io_valuReadEn_1_1;
    end
    if(when_BankedScratchMemory_l160_80) begin
      banks_0_io_reads_1_en = io_valuReadEn_1_2;
    end
    if(when_BankedScratchMemory_l160_88) begin
      banks_0_io_reads_1_en = io_valuReadEn_1_3;
    end
    if(when_BankedScratchMemory_l160_96) begin
      banks_0_io_reads_1_en = io_valuReadEn_1_4;
    end
    if(when_BankedScratchMemory_l160_104) begin
      banks_0_io_reads_1_en = io_valuReadEn_1_5;
    end
    if(when_BankedScratchMemory_l160_112) begin
      banks_0_io_reads_1_en = io_valuReadEn_1_6;
    end
    if(when_BankedScratchMemory_l160_120) begin
      banks_0_io_reads_1_en = io_valuReadEn_1_7;
    end
  end

  always @(*) begin
    banks_0_io_reads_2_addr = 8'h0;
    if(when_BankedScratchMemory_l203) begin
      if(when_BankedScratchMemory_l206) begin
        banks_0_io_reads_2_addr = scalarBankRow_0;
      end
    end
    if(when_BankedScratchMemory_l203_1) begin
      if(when_BankedScratchMemory_l206_8) begin
        banks_0_io_reads_2_addr = scalarBankRow_1;
      end
    end
    if(when_BankedScratchMemory_l203_2) begin
      if(when_BankedScratchMemory_l206_16) begin
        banks_0_io_reads_2_addr = scalarBankRow_2;
      end
    end
    if(when_BankedScratchMemory_l203_3) begin
      if(when_BankedScratchMemory_l206_24) begin
        banks_0_io_reads_2_addr = scalarBankRow_3;
      end
    end
    if(when_BankedScratchMemory_l203_4) begin
      if(when_BankedScratchMemory_l206_32) begin
        banks_0_io_reads_2_addr = scalarBankRow_4;
      end
    end
    if(when_BankedScratchMemory_l203_5) begin
      if(when_BankedScratchMemory_l206_40) begin
        banks_0_io_reads_2_addr = scalarBankRow_5;
      end
    end
    if(when_BankedScratchMemory_l203_6) begin
      if(when_BankedScratchMemory_l206_48) begin
        banks_0_io_reads_2_addr = scalarBankRow_6;
      end
    end
    if(when_BankedScratchMemory_l203_7) begin
      if(when_BankedScratchMemory_l206_56) begin
        banks_0_io_reads_2_addr = scalarBankRow_7;
      end
    end
    if(when_BankedScratchMemory_l203_8) begin
      if(when_BankedScratchMemory_l206_64) begin
        banks_0_io_reads_2_addr = scalarBankRow_8;
      end
    end
  end

  always @(*) begin
    banks_0_io_reads_2_en = 1'b0;
    if(when_BankedScratchMemory_l203) begin
      if(when_BankedScratchMemory_l206) begin
        banks_0_io_reads_2_en = 1'b1;
      end
    end
    if(when_BankedScratchMemory_l203_1) begin
      if(when_BankedScratchMemory_l206_8) begin
        banks_0_io_reads_2_en = 1'b1;
      end
    end
    if(when_BankedScratchMemory_l203_2) begin
      if(when_BankedScratchMemory_l206_16) begin
        banks_0_io_reads_2_en = 1'b1;
      end
    end
    if(when_BankedScratchMemory_l203_3) begin
      if(when_BankedScratchMemory_l206_24) begin
        banks_0_io_reads_2_en = 1'b1;
      end
    end
    if(when_BankedScratchMemory_l203_4) begin
      if(when_BankedScratchMemory_l206_32) begin
        banks_0_io_reads_2_en = 1'b1;
      end
    end
    if(when_BankedScratchMemory_l203_5) begin
      if(when_BankedScratchMemory_l206_40) begin
        banks_0_io_reads_2_en = 1'b1;
      end
    end
    if(when_BankedScratchMemory_l203_6) begin
      if(when_BankedScratchMemory_l206_48) begin
        banks_0_io_reads_2_en = 1'b1;
      end
    end
    if(when_BankedScratchMemory_l203_7) begin
      if(when_BankedScratchMemory_l206_56) begin
        banks_0_io_reads_2_en = 1'b1;
      end
    end
    if(when_BankedScratchMemory_l203_8) begin
      if(when_BankedScratchMemory_l206_64) begin
        banks_0_io_reads_2_en = 1'b1;
      end
    end
  end

  always @(*) begin
    banks_1_io_reads_0_addr = 8'h0;
    if(when_BankedScratchMemory_l160_1) begin
      banks_1_io_reads_0_addr = _zz_io_reads_0_addr;
    end
    if(when_BankedScratchMemory_l160_9) begin
      banks_1_io_reads_0_addr = _zz_io_reads_0_addr_1;
    end
    if(when_BankedScratchMemory_l160_17) begin
      banks_1_io_reads_0_addr = _zz_io_reads_0_addr_2;
    end
    if(when_BankedScratchMemory_l160_25) begin
      banks_1_io_reads_0_addr = _zz_io_reads_0_addr_3;
    end
    if(when_BankedScratchMemory_l160_33) begin
      banks_1_io_reads_0_addr = _zz_io_reads_0_addr_4;
    end
    if(when_BankedScratchMemory_l160_41) begin
      banks_1_io_reads_0_addr = _zz_io_reads_0_addr_5;
    end
    if(when_BankedScratchMemory_l160_49) begin
      banks_1_io_reads_0_addr = _zz_io_reads_0_addr_6;
    end
    if(when_BankedScratchMemory_l160_57) begin
      banks_1_io_reads_0_addr = _zz_io_reads_0_addr_7;
    end
  end

  always @(*) begin
    banks_1_io_reads_0_en = 1'b0;
    if(when_BankedScratchMemory_l160_1) begin
      banks_1_io_reads_0_en = io_valuReadEn_0_0;
    end
    if(when_BankedScratchMemory_l160_9) begin
      banks_1_io_reads_0_en = io_valuReadEn_0_1;
    end
    if(when_BankedScratchMemory_l160_17) begin
      banks_1_io_reads_0_en = io_valuReadEn_0_2;
    end
    if(when_BankedScratchMemory_l160_25) begin
      banks_1_io_reads_0_en = io_valuReadEn_0_3;
    end
    if(when_BankedScratchMemory_l160_33) begin
      banks_1_io_reads_0_en = io_valuReadEn_0_4;
    end
    if(when_BankedScratchMemory_l160_41) begin
      banks_1_io_reads_0_en = io_valuReadEn_0_5;
    end
    if(when_BankedScratchMemory_l160_49) begin
      banks_1_io_reads_0_en = io_valuReadEn_0_6;
    end
    if(when_BankedScratchMemory_l160_57) begin
      banks_1_io_reads_0_en = io_valuReadEn_0_7;
    end
  end

  always @(*) begin
    banks_1_io_reads_1_addr = 8'h0;
    if(when_BankedScratchMemory_l160_65) begin
      banks_1_io_reads_1_addr = _zz_io_reads_1_addr;
    end
    if(when_BankedScratchMemory_l160_73) begin
      banks_1_io_reads_1_addr = _zz_io_reads_1_addr_1;
    end
    if(when_BankedScratchMemory_l160_81) begin
      banks_1_io_reads_1_addr = _zz_io_reads_1_addr_2;
    end
    if(when_BankedScratchMemory_l160_89) begin
      banks_1_io_reads_1_addr = _zz_io_reads_1_addr_3;
    end
    if(when_BankedScratchMemory_l160_97) begin
      banks_1_io_reads_1_addr = _zz_io_reads_1_addr_4;
    end
    if(when_BankedScratchMemory_l160_105) begin
      banks_1_io_reads_1_addr = _zz_io_reads_1_addr_5;
    end
    if(when_BankedScratchMemory_l160_113) begin
      banks_1_io_reads_1_addr = _zz_io_reads_1_addr_6;
    end
    if(when_BankedScratchMemory_l160_121) begin
      banks_1_io_reads_1_addr = _zz_io_reads_1_addr_7;
    end
  end

  always @(*) begin
    banks_1_io_reads_1_en = 1'b0;
    if(when_BankedScratchMemory_l160_65) begin
      banks_1_io_reads_1_en = io_valuReadEn_1_0;
    end
    if(when_BankedScratchMemory_l160_73) begin
      banks_1_io_reads_1_en = io_valuReadEn_1_1;
    end
    if(when_BankedScratchMemory_l160_81) begin
      banks_1_io_reads_1_en = io_valuReadEn_1_2;
    end
    if(when_BankedScratchMemory_l160_89) begin
      banks_1_io_reads_1_en = io_valuReadEn_1_3;
    end
    if(when_BankedScratchMemory_l160_97) begin
      banks_1_io_reads_1_en = io_valuReadEn_1_4;
    end
    if(when_BankedScratchMemory_l160_105) begin
      banks_1_io_reads_1_en = io_valuReadEn_1_5;
    end
    if(when_BankedScratchMemory_l160_113) begin
      banks_1_io_reads_1_en = io_valuReadEn_1_6;
    end
    if(when_BankedScratchMemory_l160_121) begin
      banks_1_io_reads_1_en = io_valuReadEn_1_7;
    end
  end

  always @(*) begin
    banks_1_io_reads_2_addr = 8'h0;
    if(when_BankedScratchMemory_l203) begin
      if(when_BankedScratchMemory_l206_1) begin
        banks_1_io_reads_2_addr = scalarBankRow_0;
      end
    end
    if(when_BankedScratchMemory_l203_1) begin
      if(when_BankedScratchMemory_l206_9) begin
        banks_1_io_reads_2_addr = scalarBankRow_1;
      end
    end
    if(when_BankedScratchMemory_l203_2) begin
      if(when_BankedScratchMemory_l206_17) begin
        banks_1_io_reads_2_addr = scalarBankRow_2;
      end
    end
    if(when_BankedScratchMemory_l203_3) begin
      if(when_BankedScratchMemory_l206_25) begin
        banks_1_io_reads_2_addr = scalarBankRow_3;
      end
    end
    if(when_BankedScratchMemory_l203_4) begin
      if(when_BankedScratchMemory_l206_33) begin
        banks_1_io_reads_2_addr = scalarBankRow_4;
      end
    end
    if(when_BankedScratchMemory_l203_5) begin
      if(when_BankedScratchMemory_l206_41) begin
        banks_1_io_reads_2_addr = scalarBankRow_5;
      end
    end
    if(when_BankedScratchMemory_l203_6) begin
      if(when_BankedScratchMemory_l206_49) begin
        banks_1_io_reads_2_addr = scalarBankRow_6;
      end
    end
    if(when_BankedScratchMemory_l203_7) begin
      if(when_BankedScratchMemory_l206_57) begin
        banks_1_io_reads_2_addr = scalarBankRow_7;
      end
    end
    if(when_BankedScratchMemory_l203_8) begin
      if(when_BankedScratchMemory_l206_65) begin
        banks_1_io_reads_2_addr = scalarBankRow_8;
      end
    end
  end

  always @(*) begin
    banks_1_io_reads_2_en = 1'b0;
    if(when_BankedScratchMemory_l203) begin
      if(when_BankedScratchMemory_l206_1) begin
        banks_1_io_reads_2_en = 1'b1;
      end
    end
    if(when_BankedScratchMemory_l203_1) begin
      if(when_BankedScratchMemory_l206_9) begin
        banks_1_io_reads_2_en = 1'b1;
      end
    end
    if(when_BankedScratchMemory_l203_2) begin
      if(when_BankedScratchMemory_l206_17) begin
        banks_1_io_reads_2_en = 1'b1;
      end
    end
    if(when_BankedScratchMemory_l203_3) begin
      if(when_BankedScratchMemory_l206_25) begin
        banks_1_io_reads_2_en = 1'b1;
      end
    end
    if(when_BankedScratchMemory_l203_4) begin
      if(when_BankedScratchMemory_l206_33) begin
        banks_1_io_reads_2_en = 1'b1;
      end
    end
    if(when_BankedScratchMemory_l203_5) begin
      if(when_BankedScratchMemory_l206_41) begin
        banks_1_io_reads_2_en = 1'b1;
      end
    end
    if(when_BankedScratchMemory_l203_6) begin
      if(when_BankedScratchMemory_l206_49) begin
        banks_1_io_reads_2_en = 1'b1;
      end
    end
    if(when_BankedScratchMemory_l203_7) begin
      if(when_BankedScratchMemory_l206_57) begin
        banks_1_io_reads_2_en = 1'b1;
      end
    end
    if(when_BankedScratchMemory_l203_8) begin
      if(when_BankedScratchMemory_l206_65) begin
        banks_1_io_reads_2_en = 1'b1;
      end
    end
  end

  always @(*) begin
    banks_2_io_reads_0_addr = 8'h0;
    if(when_BankedScratchMemory_l160_2) begin
      banks_2_io_reads_0_addr = _zz_io_reads_0_addr;
    end
    if(when_BankedScratchMemory_l160_10) begin
      banks_2_io_reads_0_addr = _zz_io_reads_0_addr_1;
    end
    if(when_BankedScratchMemory_l160_18) begin
      banks_2_io_reads_0_addr = _zz_io_reads_0_addr_2;
    end
    if(when_BankedScratchMemory_l160_26) begin
      banks_2_io_reads_0_addr = _zz_io_reads_0_addr_3;
    end
    if(when_BankedScratchMemory_l160_34) begin
      banks_2_io_reads_0_addr = _zz_io_reads_0_addr_4;
    end
    if(when_BankedScratchMemory_l160_42) begin
      banks_2_io_reads_0_addr = _zz_io_reads_0_addr_5;
    end
    if(when_BankedScratchMemory_l160_50) begin
      banks_2_io_reads_0_addr = _zz_io_reads_0_addr_6;
    end
    if(when_BankedScratchMemory_l160_58) begin
      banks_2_io_reads_0_addr = _zz_io_reads_0_addr_7;
    end
  end

  always @(*) begin
    banks_2_io_reads_0_en = 1'b0;
    if(when_BankedScratchMemory_l160_2) begin
      banks_2_io_reads_0_en = io_valuReadEn_0_0;
    end
    if(when_BankedScratchMemory_l160_10) begin
      banks_2_io_reads_0_en = io_valuReadEn_0_1;
    end
    if(when_BankedScratchMemory_l160_18) begin
      banks_2_io_reads_0_en = io_valuReadEn_0_2;
    end
    if(when_BankedScratchMemory_l160_26) begin
      banks_2_io_reads_0_en = io_valuReadEn_0_3;
    end
    if(when_BankedScratchMemory_l160_34) begin
      banks_2_io_reads_0_en = io_valuReadEn_0_4;
    end
    if(when_BankedScratchMemory_l160_42) begin
      banks_2_io_reads_0_en = io_valuReadEn_0_5;
    end
    if(when_BankedScratchMemory_l160_50) begin
      banks_2_io_reads_0_en = io_valuReadEn_0_6;
    end
    if(when_BankedScratchMemory_l160_58) begin
      banks_2_io_reads_0_en = io_valuReadEn_0_7;
    end
  end

  always @(*) begin
    banks_2_io_reads_1_addr = 8'h0;
    if(when_BankedScratchMemory_l160_66) begin
      banks_2_io_reads_1_addr = _zz_io_reads_1_addr;
    end
    if(when_BankedScratchMemory_l160_74) begin
      banks_2_io_reads_1_addr = _zz_io_reads_1_addr_1;
    end
    if(when_BankedScratchMemory_l160_82) begin
      banks_2_io_reads_1_addr = _zz_io_reads_1_addr_2;
    end
    if(when_BankedScratchMemory_l160_90) begin
      banks_2_io_reads_1_addr = _zz_io_reads_1_addr_3;
    end
    if(when_BankedScratchMemory_l160_98) begin
      banks_2_io_reads_1_addr = _zz_io_reads_1_addr_4;
    end
    if(when_BankedScratchMemory_l160_106) begin
      banks_2_io_reads_1_addr = _zz_io_reads_1_addr_5;
    end
    if(when_BankedScratchMemory_l160_114) begin
      banks_2_io_reads_1_addr = _zz_io_reads_1_addr_6;
    end
    if(when_BankedScratchMemory_l160_122) begin
      banks_2_io_reads_1_addr = _zz_io_reads_1_addr_7;
    end
  end

  always @(*) begin
    banks_2_io_reads_1_en = 1'b0;
    if(when_BankedScratchMemory_l160_66) begin
      banks_2_io_reads_1_en = io_valuReadEn_1_0;
    end
    if(when_BankedScratchMemory_l160_74) begin
      banks_2_io_reads_1_en = io_valuReadEn_1_1;
    end
    if(when_BankedScratchMemory_l160_82) begin
      banks_2_io_reads_1_en = io_valuReadEn_1_2;
    end
    if(when_BankedScratchMemory_l160_90) begin
      banks_2_io_reads_1_en = io_valuReadEn_1_3;
    end
    if(when_BankedScratchMemory_l160_98) begin
      banks_2_io_reads_1_en = io_valuReadEn_1_4;
    end
    if(when_BankedScratchMemory_l160_106) begin
      banks_2_io_reads_1_en = io_valuReadEn_1_5;
    end
    if(when_BankedScratchMemory_l160_114) begin
      banks_2_io_reads_1_en = io_valuReadEn_1_6;
    end
    if(when_BankedScratchMemory_l160_122) begin
      banks_2_io_reads_1_en = io_valuReadEn_1_7;
    end
  end

  always @(*) begin
    banks_2_io_reads_2_addr = 8'h0;
    if(when_BankedScratchMemory_l203) begin
      if(when_BankedScratchMemory_l206_2) begin
        banks_2_io_reads_2_addr = scalarBankRow_0;
      end
    end
    if(when_BankedScratchMemory_l203_1) begin
      if(when_BankedScratchMemory_l206_10) begin
        banks_2_io_reads_2_addr = scalarBankRow_1;
      end
    end
    if(when_BankedScratchMemory_l203_2) begin
      if(when_BankedScratchMemory_l206_18) begin
        banks_2_io_reads_2_addr = scalarBankRow_2;
      end
    end
    if(when_BankedScratchMemory_l203_3) begin
      if(when_BankedScratchMemory_l206_26) begin
        banks_2_io_reads_2_addr = scalarBankRow_3;
      end
    end
    if(when_BankedScratchMemory_l203_4) begin
      if(when_BankedScratchMemory_l206_34) begin
        banks_2_io_reads_2_addr = scalarBankRow_4;
      end
    end
    if(when_BankedScratchMemory_l203_5) begin
      if(when_BankedScratchMemory_l206_42) begin
        banks_2_io_reads_2_addr = scalarBankRow_5;
      end
    end
    if(when_BankedScratchMemory_l203_6) begin
      if(when_BankedScratchMemory_l206_50) begin
        banks_2_io_reads_2_addr = scalarBankRow_6;
      end
    end
    if(when_BankedScratchMemory_l203_7) begin
      if(when_BankedScratchMemory_l206_58) begin
        banks_2_io_reads_2_addr = scalarBankRow_7;
      end
    end
    if(when_BankedScratchMemory_l203_8) begin
      if(when_BankedScratchMemory_l206_66) begin
        banks_2_io_reads_2_addr = scalarBankRow_8;
      end
    end
  end

  always @(*) begin
    banks_2_io_reads_2_en = 1'b0;
    if(when_BankedScratchMemory_l203) begin
      if(when_BankedScratchMemory_l206_2) begin
        banks_2_io_reads_2_en = 1'b1;
      end
    end
    if(when_BankedScratchMemory_l203_1) begin
      if(when_BankedScratchMemory_l206_10) begin
        banks_2_io_reads_2_en = 1'b1;
      end
    end
    if(when_BankedScratchMemory_l203_2) begin
      if(when_BankedScratchMemory_l206_18) begin
        banks_2_io_reads_2_en = 1'b1;
      end
    end
    if(when_BankedScratchMemory_l203_3) begin
      if(when_BankedScratchMemory_l206_26) begin
        banks_2_io_reads_2_en = 1'b1;
      end
    end
    if(when_BankedScratchMemory_l203_4) begin
      if(when_BankedScratchMemory_l206_34) begin
        banks_2_io_reads_2_en = 1'b1;
      end
    end
    if(when_BankedScratchMemory_l203_5) begin
      if(when_BankedScratchMemory_l206_42) begin
        banks_2_io_reads_2_en = 1'b1;
      end
    end
    if(when_BankedScratchMemory_l203_6) begin
      if(when_BankedScratchMemory_l206_50) begin
        banks_2_io_reads_2_en = 1'b1;
      end
    end
    if(when_BankedScratchMemory_l203_7) begin
      if(when_BankedScratchMemory_l206_58) begin
        banks_2_io_reads_2_en = 1'b1;
      end
    end
    if(when_BankedScratchMemory_l203_8) begin
      if(when_BankedScratchMemory_l206_66) begin
        banks_2_io_reads_2_en = 1'b1;
      end
    end
  end

  always @(*) begin
    banks_3_io_reads_0_addr = 8'h0;
    if(when_BankedScratchMemory_l160_3) begin
      banks_3_io_reads_0_addr = _zz_io_reads_0_addr;
    end
    if(when_BankedScratchMemory_l160_11) begin
      banks_3_io_reads_0_addr = _zz_io_reads_0_addr_1;
    end
    if(when_BankedScratchMemory_l160_19) begin
      banks_3_io_reads_0_addr = _zz_io_reads_0_addr_2;
    end
    if(when_BankedScratchMemory_l160_27) begin
      banks_3_io_reads_0_addr = _zz_io_reads_0_addr_3;
    end
    if(when_BankedScratchMemory_l160_35) begin
      banks_3_io_reads_0_addr = _zz_io_reads_0_addr_4;
    end
    if(when_BankedScratchMemory_l160_43) begin
      banks_3_io_reads_0_addr = _zz_io_reads_0_addr_5;
    end
    if(when_BankedScratchMemory_l160_51) begin
      banks_3_io_reads_0_addr = _zz_io_reads_0_addr_6;
    end
    if(when_BankedScratchMemory_l160_59) begin
      banks_3_io_reads_0_addr = _zz_io_reads_0_addr_7;
    end
  end

  always @(*) begin
    banks_3_io_reads_0_en = 1'b0;
    if(when_BankedScratchMemory_l160_3) begin
      banks_3_io_reads_0_en = io_valuReadEn_0_0;
    end
    if(when_BankedScratchMemory_l160_11) begin
      banks_3_io_reads_0_en = io_valuReadEn_0_1;
    end
    if(when_BankedScratchMemory_l160_19) begin
      banks_3_io_reads_0_en = io_valuReadEn_0_2;
    end
    if(when_BankedScratchMemory_l160_27) begin
      banks_3_io_reads_0_en = io_valuReadEn_0_3;
    end
    if(when_BankedScratchMemory_l160_35) begin
      banks_3_io_reads_0_en = io_valuReadEn_0_4;
    end
    if(when_BankedScratchMemory_l160_43) begin
      banks_3_io_reads_0_en = io_valuReadEn_0_5;
    end
    if(when_BankedScratchMemory_l160_51) begin
      banks_3_io_reads_0_en = io_valuReadEn_0_6;
    end
    if(when_BankedScratchMemory_l160_59) begin
      banks_3_io_reads_0_en = io_valuReadEn_0_7;
    end
  end

  always @(*) begin
    banks_3_io_reads_1_addr = 8'h0;
    if(when_BankedScratchMemory_l160_67) begin
      banks_3_io_reads_1_addr = _zz_io_reads_1_addr;
    end
    if(when_BankedScratchMemory_l160_75) begin
      banks_3_io_reads_1_addr = _zz_io_reads_1_addr_1;
    end
    if(when_BankedScratchMemory_l160_83) begin
      banks_3_io_reads_1_addr = _zz_io_reads_1_addr_2;
    end
    if(when_BankedScratchMemory_l160_91) begin
      banks_3_io_reads_1_addr = _zz_io_reads_1_addr_3;
    end
    if(when_BankedScratchMemory_l160_99) begin
      banks_3_io_reads_1_addr = _zz_io_reads_1_addr_4;
    end
    if(when_BankedScratchMemory_l160_107) begin
      banks_3_io_reads_1_addr = _zz_io_reads_1_addr_5;
    end
    if(when_BankedScratchMemory_l160_115) begin
      banks_3_io_reads_1_addr = _zz_io_reads_1_addr_6;
    end
    if(when_BankedScratchMemory_l160_123) begin
      banks_3_io_reads_1_addr = _zz_io_reads_1_addr_7;
    end
  end

  always @(*) begin
    banks_3_io_reads_1_en = 1'b0;
    if(when_BankedScratchMemory_l160_67) begin
      banks_3_io_reads_1_en = io_valuReadEn_1_0;
    end
    if(when_BankedScratchMemory_l160_75) begin
      banks_3_io_reads_1_en = io_valuReadEn_1_1;
    end
    if(when_BankedScratchMemory_l160_83) begin
      banks_3_io_reads_1_en = io_valuReadEn_1_2;
    end
    if(when_BankedScratchMemory_l160_91) begin
      banks_3_io_reads_1_en = io_valuReadEn_1_3;
    end
    if(when_BankedScratchMemory_l160_99) begin
      banks_3_io_reads_1_en = io_valuReadEn_1_4;
    end
    if(when_BankedScratchMemory_l160_107) begin
      banks_3_io_reads_1_en = io_valuReadEn_1_5;
    end
    if(when_BankedScratchMemory_l160_115) begin
      banks_3_io_reads_1_en = io_valuReadEn_1_6;
    end
    if(when_BankedScratchMemory_l160_123) begin
      banks_3_io_reads_1_en = io_valuReadEn_1_7;
    end
  end

  always @(*) begin
    banks_3_io_reads_2_addr = 8'h0;
    if(when_BankedScratchMemory_l203) begin
      if(when_BankedScratchMemory_l206_3) begin
        banks_3_io_reads_2_addr = scalarBankRow_0;
      end
    end
    if(when_BankedScratchMemory_l203_1) begin
      if(when_BankedScratchMemory_l206_11) begin
        banks_3_io_reads_2_addr = scalarBankRow_1;
      end
    end
    if(when_BankedScratchMemory_l203_2) begin
      if(when_BankedScratchMemory_l206_19) begin
        banks_3_io_reads_2_addr = scalarBankRow_2;
      end
    end
    if(when_BankedScratchMemory_l203_3) begin
      if(when_BankedScratchMemory_l206_27) begin
        banks_3_io_reads_2_addr = scalarBankRow_3;
      end
    end
    if(when_BankedScratchMemory_l203_4) begin
      if(when_BankedScratchMemory_l206_35) begin
        banks_3_io_reads_2_addr = scalarBankRow_4;
      end
    end
    if(when_BankedScratchMemory_l203_5) begin
      if(when_BankedScratchMemory_l206_43) begin
        banks_3_io_reads_2_addr = scalarBankRow_5;
      end
    end
    if(when_BankedScratchMemory_l203_6) begin
      if(when_BankedScratchMemory_l206_51) begin
        banks_3_io_reads_2_addr = scalarBankRow_6;
      end
    end
    if(when_BankedScratchMemory_l203_7) begin
      if(when_BankedScratchMemory_l206_59) begin
        banks_3_io_reads_2_addr = scalarBankRow_7;
      end
    end
    if(when_BankedScratchMemory_l203_8) begin
      if(when_BankedScratchMemory_l206_67) begin
        banks_3_io_reads_2_addr = scalarBankRow_8;
      end
    end
  end

  always @(*) begin
    banks_3_io_reads_2_en = 1'b0;
    if(when_BankedScratchMemory_l203) begin
      if(when_BankedScratchMemory_l206_3) begin
        banks_3_io_reads_2_en = 1'b1;
      end
    end
    if(when_BankedScratchMemory_l203_1) begin
      if(when_BankedScratchMemory_l206_11) begin
        banks_3_io_reads_2_en = 1'b1;
      end
    end
    if(when_BankedScratchMemory_l203_2) begin
      if(when_BankedScratchMemory_l206_19) begin
        banks_3_io_reads_2_en = 1'b1;
      end
    end
    if(when_BankedScratchMemory_l203_3) begin
      if(when_BankedScratchMemory_l206_27) begin
        banks_3_io_reads_2_en = 1'b1;
      end
    end
    if(when_BankedScratchMemory_l203_4) begin
      if(when_BankedScratchMemory_l206_35) begin
        banks_3_io_reads_2_en = 1'b1;
      end
    end
    if(when_BankedScratchMemory_l203_5) begin
      if(when_BankedScratchMemory_l206_43) begin
        banks_3_io_reads_2_en = 1'b1;
      end
    end
    if(when_BankedScratchMemory_l203_6) begin
      if(when_BankedScratchMemory_l206_51) begin
        banks_3_io_reads_2_en = 1'b1;
      end
    end
    if(when_BankedScratchMemory_l203_7) begin
      if(when_BankedScratchMemory_l206_59) begin
        banks_3_io_reads_2_en = 1'b1;
      end
    end
    if(when_BankedScratchMemory_l203_8) begin
      if(when_BankedScratchMemory_l206_67) begin
        banks_3_io_reads_2_en = 1'b1;
      end
    end
  end

  always @(*) begin
    banks_4_io_reads_0_addr = 8'h0;
    if(when_BankedScratchMemory_l160_4) begin
      banks_4_io_reads_0_addr = _zz_io_reads_0_addr;
    end
    if(when_BankedScratchMemory_l160_12) begin
      banks_4_io_reads_0_addr = _zz_io_reads_0_addr_1;
    end
    if(when_BankedScratchMemory_l160_20) begin
      banks_4_io_reads_0_addr = _zz_io_reads_0_addr_2;
    end
    if(when_BankedScratchMemory_l160_28) begin
      banks_4_io_reads_0_addr = _zz_io_reads_0_addr_3;
    end
    if(when_BankedScratchMemory_l160_36) begin
      banks_4_io_reads_0_addr = _zz_io_reads_0_addr_4;
    end
    if(when_BankedScratchMemory_l160_44) begin
      banks_4_io_reads_0_addr = _zz_io_reads_0_addr_5;
    end
    if(when_BankedScratchMemory_l160_52) begin
      banks_4_io_reads_0_addr = _zz_io_reads_0_addr_6;
    end
    if(when_BankedScratchMemory_l160_60) begin
      banks_4_io_reads_0_addr = _zz_io_reads_0_addr_7;
    end
  end

  always @(*) begin
    banks_4_io_reads_0_en = 1'b0;
    if(when_BankedScratchMemory_l160_4) begin
      banks_4_io_reads_0_en = io_valuReadEn_0_0;
    end
    if(when_BankedScratchMemory_l160_12) begin
      banks_4_io_reads_0_en = io_valuReadEn_0_1;
    end
    if(when_BankedScratchMemory_l160_20) begin
      banks_4_io_reads_0_en = io_valuReadEn_0_2;
    end
    if(when_BankedScratchMemory_l160_28) begin
      banks_4_io_reads_0_en = io_valuReadEn_0_3;
    end
    if(when_BankedScratchMemory_l160_36) begin
      banks_4_io_reads_0_en = io_valuReadEn_0_4;
    end
    if(when_BankedScratchMemory_l160_44) begin
      banks_4_io_reads_0_en = io_valuReadEn_0_5;
    end
    if(when_BankedScratchMemory_l160_52) begin
      banks_4_io_reads_0_en = io_valuReadEn_0_6;
    end
    if(when_BankedScratchMemory_l160_60) begin
      banks_4_io_reads_0_en = io_valuReadEn_0_7;
    end
  end

  always @(*) begin
    banks_4_io_reads_1_addr = 8'h0;
    if(when_BankedScratchMemory_l160_68) begin
      banks_4_io_reads_1_addr = _zz_io_reads_1_addr;
    end
    if(when_BankedScratchMemory_l160_76) begin
      banks_4_io_reads_1_addr = _zz_io_reads_1_addr_1;
    end
    if(when_BankedScratchMemory_l160_84) begin
      banks_4_io_reads_1_addr = _zz_io_reads_1_addr_2;
    end
    if(when_BankedScratchMemory_l160_92) begin
      banks_4_io_reads_1_addr = _zz_io_reads_1_addr_3;
    end
    if(when_BankedScratchMemory_l160_100) begin
      banks_4_io_reads_1_addr = _zz_io_reads_1_addr_4;
    end
    if(when_BankedScratchMemory_l160_108) begin
      banks_4_io_reads_1_addr = _zz_io_reads_1_addr_5;
    end
    if(when_BankedScratchMemory_l160_116) begin
      banks_4_io_reads_1_addr = _zz_io_reads_1_addr_6;
    end
    if(when_BankedScratchMemory_l160_124) begin
      banks_4_io_reads_1_addr = _zz_io_reads_1_addr_7;
    end
  end

  always @(*) begin
    banks_4_io_reads_1_en = 1'b0;
    if(when_BankedScratchMemory_l160_68) begin
      banks_4_io_reads_1_en = io_valuReadEn_1_0;
    end
    if(when_BankedScratchMemory_l160_76) begin
      banks_4_io_reads_1_en = io_valuReadEn_1_1;
    end
    if(when_BankedScratchMemory_l160_84) begin
      banks_4_io_reads_1_en = io_valuReadEn_1_2;
    end
    if(when_BankedScratchMemory_l160_92) begin
      banks_4_io_reads_1_en = io_valuReadEn_1_3;
    end
    if(when_BankedScratchMemory_l160_100) begin
      banks_4_io_reads_1_en = io_valuReadEn_1_4;
    end
    if(when_BankedScratchMemory_l160_108) begin
      banks_4_io_reads_1_en = io_valuReadEn_1_5;
    end
    if(when_BankedScratchMemory_l160_116) begin
      banks_4_io_reads_1_en = io_valuReadEn_1_6;
    end
    if(when_BankedScratchMemory_l160_124) begin
      banks_4_io_reads_1_en = io_valuReadEn_1_7;
    end
  end

  always @(*) begin
    banks_4_io_reads_2_addr = 8'h0;
    if(when_BankedScratchMemory_l203) begin
      if(when_BankedScratchMemory_l206_4) begin
        banks_4_io_reads_2_addr = scalarBankRow_0;
      end
    end
    if(when_BankedScratchMemory_l203_1) begin
      if(when_BankedScratchMemory_l206_12) begin
        banks_4_io_reads_2_addr = scalarBankRow_1;
      end
    end
    if(when_BankedScratchMemory_l203_2) begin
      if(when_BankedScratchMemory_l206_20) begin
        banks_4_io_reads_2_addr = scalarBankRow_2;
      end
    end
    if(when_BankedScratchMemory_l203_3) begin
      if(when_BankedScratchMemory_l206_28) begin
        banks_4_io_reads_2_addr = scalarBankRow_3;
      end
    end
    if(when_BankedScratchMemory_l203_4) begin
      if(when_BankedScratchMemory_l206_36) begin
        banks_4_io_reads_2_addr = scalarBankRow_4;
      end
    end
    if(when_BankedScratchMemory_l203_5) begin
      if(when_BankedScratchMemory_l206_44) begin
        banks_4_io_reads_2_addr = scalarBankRow_5;
      end
    end
    if(when_BankedScratchMemory_l203_6) begin
      if(when_BankedScratchMemory_l206_52) begin
        banks_4_io_reads_2_addr = scalarBankRow_6;
      end
    end
    if(when_BankedScratchMemory_l203_7) begin
      if(when_BankedScratchMemory_l206_60) begin
        banks_4_io_reads_2_addr = scalarBankRow_7;
      end
    end
    if(when_BankedScratchMemory_l203_8) begin
      if(when_BankedScratchMemory_l206_68) begin
        banks_4_io_reads_2_addr = scalarBankRow_8;
      end
    end
  end

  always @(*) begin
    banks_4_io_reads_2_en = 1'b0;
    if(when_BankedScratchMemory_l203) begin
      if(when_BankedScratchMemory_l206_4) begin
        banks_4_io_reads_2_en = 1'b1;
      end
    end
    if(when_BankedScratchMemory_l203_1) begin
      if(when_BankedScratchMemory_l206_12) begin
        banks_4_io_reads_2_en = 1'b1;
      end
    end
    if(when_BankedScratchMemory_l203_2) begin
      if(when_BankedScratchMemory_l206_20) begin
        banks_4_io_reads_2_en = 1'b1;
      end
    end
    if(when_BankedScratchMemory_l203_3) begin
      if(when_BankedScratchMemory_l206_28) begin
        banks_4_io_reads_2_en = 1'b1;
      end
    end
    if(when_BankedScratchMemory_l203_4) begin
      if(when_BankedScratchMemory_l206_36) begin
        banks_4_io_reads_2_en = 1'b1;
      end
    end
    if(when_BankedScratchMemory_l203_5) begin
      if(when_BankedScratchMemory_l206_44) begin
        banks_4_io_reads_2_en = 1'b1;
      end
    end
    if(when_BankedScratchMemory_l203_6) begin
      if(when_BankedScratchMemory_l206_52) begin
        banks_4_io_reads_2_en = 1'b1;
      end
    end
    if(when_BankedScratchMemory_l203_7) begin
      if(when_BankedScratchMemory_l206_60) begin
        banks_4_io_reads_2_en = 1'b1;
      end
    end
    if(when_BankedScratchMemory_l203_8) begin
      if(when_BankedScratchMemory_l206_68) begin
        banks_4_io_reads_2_en = 1'b1;
      end
    end
  end

  always @(*) begin
    banks_5_io_reads_0_addr = 8'h0;
    if(when_BankedScratchMemory_l160_5) begin
      banks_5_io_reads_0_addr = _zz_io_reads_0_addr;
    end
    if(when_BankedScratchMemory_l160_13) begin
      banks_5_io_reads_0_addr = _zz_io_reads_0_addr_1;
    end
    if(when_BankedScratchMemory_l160_21) begin
      banks_5_io_reads_0_addr = _zz_io_reads_0_addr_2;
    end
    if(when_BankedScratchMemory_l160_29) begin
      banks_5_io_reads_0_addr = _zz_io_reads_0_addr_3;
    end
    if(when_BankedScratchMemory_l160_37) begin
      banks_5_io_reads_0_addr = _zz_io_reads_0_addr_4;
    end
    if(when_BankedScratchMemory_l160_45) begin
      banks_5_io_reads_0_addr = _zz_io_reads_0_addr_5;
    end
    if(when_BankedScratchMemory_l160_53) begin
      banks_5_io_reads_0_addr = _zz_io_reads_0_addr_6;
    end
    if(when_BankedScratchMemory_l160_61) begin
      banks_5_io_reads_0_addr = _zz_io_reads_0_addr_7;
    end
  end

  always @(*) begin
    banks_5_io_reads_0_en = 1'b0;
    if(when_BankedScratchMemory_l160_5) begin
      banks_5_io_reads_0_en = io_valuReadEn_0_0;
    end
    if(when_BankedScratchMemory_l160_13) begin
      banks_5_io_reads_0_en = io_valuReadEn_0_1;
    end
    if(when_BankedScratchMemory_l160_21) begin
      banks_5_io_reads_0_en = io_valuReadEn_0_2;
    end
    if(when_BankedScratchMemory_l160_29) begin
      banks_5_io_reads_0_en = io_valuReadEn_0_3;
    end
    if(when_BankedScratchMemory_l160_37) begin
      banks_5_io_reads_0_en = io_valuReadEn_0_4;
    end
    if(when_BankedScratchMemory_l160_45) begin
      banks_5_io_reads_0_en = io_valuReadEn_0_5;
    end
    if(when_BankedScratchMemory_l160_53) begin
      banks_5_io_reads_0_en = io_valuReadEn_0_6;
    end
    if(when_BankedScratchMemory_l160_61) begin
      banks_5_io_reads_0_en = io_valuReadEn_0_7;
    end
  end

  always @(*) begin
    banks_5_io_reads_1_addr = 8'h0;
    if(when_BankedScratchMemory_l160_69) begin
      banks_5_io_reads_1_addr = _zz_io_reads_1_addr;
    end
    if(when_BankedScratchMemory_l160_77) begin
      banks_5_io_reads_1_addr = _zz_io_reads_1_addr_1;
    end
    if(when_BankedScratchMemory_l160_85) begin
      banks_5_io_reads_1_addr = _zz_io_reads_1_addr_2;
    end
    if(when_BankedScratchMemory_l160_93) begin
      banks_5_io_reads_1_addr = _zz_io_reads_1_addr_3;
    end
    if(when_BankedScratchMemory_l160_101) begin
      banks_5_io_reads_1_addr = _zz_io_reads_1_addr_4;
    end
    if(when_BankedScratchMemory_l160_109) begin
      banks_5_io_reads_1_addr = _zz_io_reads_1_addr_5;
    end
    if(when_BankedScratchMemory_l160_117) begin
      banks_5_io_reads_1_addr = _zz_io_reads_1_addr_6;
    end
    if(when_BankedScratchMemory_l160_125) begin
      banks_5_io_reads_1_addr = _zz_io_reads_1_addr_7;
    end
  end

  always @(*) begin
    banks_5_io_reads_1_en = 1'b0;
    if(when_BankedScratchMemory_l160_69) begin
      banks_5_io_reads_1_en = io_valuReadEn_1_0;
    end
    if(when_BankedScratchMemory_l160_77) begin
      banks_5_io_reads_1_en = io_valuReadEn_1_1;
    end
    if(when_BankedScratchMemory_l160_85) begin
      banks_5_io_reads_1_en = io_valuReadEn_1_2;
    end
    if(when_BankedScratchMemory_l160_93) begin
      banks_5_io_reads_1_en = io_valuReadEn_1_3;
    end
    if(when_BankedScratchMemory_l160_101) begin
      banks_5_io_reads_1_en = io_valuReadEn_1_4;
    end
    if(when_BankedScratchMemory_l160_109) begin
      banks_5_io_reads_1_en = io_valuReadEn_1_5;
    end
    if(when_BankedScratchMemory_l160_117) begin
      banks_5_io_reads_1_en = io_valuReadEn_1_6;
    end
    if(when_BankedScratchMemory_l160_125) begin
      banks_5_io_reads_1_en = io_valuReadEn_1_7;
    end
  end

  always @(*) begin
    banks_5_io_reads_2_addr = 8'h0;
    if(when_BankedScratchMemory_l203) begin
      if(when_BankedScratchMemory_l206_5) begin
        banks_5_io_reads_2_addr = scalarBankRow_0;
      end
    end
    if(when_BankedScratchMemory_l203_1) begin
      if(when_BankedScratchMemory_l206_13) begin
        banks_5_io_reads_2_addr = scalarBankRow_1;
      end
    end
    if(when_BankedScratchMemory_l203_2) begin
      if(when_BankedScratchMemory_l206_21) begin
        banks_5_io_reads_2_addr = scalarBankRow_2;
      end
    end
    if(when_BankedScratchMemory_l203_3) begin
      if(when_BankedScratchMemory_l206_29) begin
        banks_5_io_reads_2_addr = scalarBankRow_3;
      end
    end
    if(when_BankedScratchMemory_l203_4) begin
      if(when_BankedScratchMemory_l206_37) begin
        banks_5_io_reads_2_addr = scalarBankRow_4;
      end
    end
    if(when_BankedScratchMemory_l203_5) begin
      if(when_BankedScratchMemory_l206_45) begin
        banks_5_io_reads_2_addr = scalarBankRow_5;
      end
    end
    if(when_BankedScratchMemory_l203_6) begin
      if(when_BankedScratchMemory_l206_53) begin
        banks_5_io_reads_2_addr = scalarBankRow_6;
      end
    end
    if(when_BankedScratchMemory_l203_7) begin
      if(when_BankedScratchMemory_l206_61) begin
        banks_5_io_reads_2_addr = scalarBankRow_7;
      end
    end
    if(when_BankedScratchMemory_l203_8) begin
      if(when_BankedScratchMemory_l206_69) begin
        banks_5_io_reads_2_addr = scalarBankRow_8;
      end
    end
  end

  always @(*) begin
    banks_5_io_reads_2_en = 1'b0;
    if(when_BankedScratchMemory_l203) begin
      if(when_BankedScratchMemory_l206_5) begin
        banks_5_io_reads_2_en = 1'b1;
      end
    end
    if(when_BankedScratchMemory_l203_1) begin
      if(when_BankedScratchMemory_l206_13) begin
        banks_5_io_reads_2_en = 1'b1;
      end
    end
    if(when_BankedScratchMemory_l203_2) begin
      if(when_BankedScratchMemory_l206_21) begin
        banks_5_io_reads_2_en = 1'b1;
      end
    end
    if(when_BankedScratchMemory_l203_3) begin
      if(when_BankedScratchMemory_l206_29) begin
        banks_5_io_reads_2_en = 1'b1;
      end
    end
    if(when_BankedScratchMemory_l203_4) begin
      if(when_BankedScratchMemory_l206_37) begin
        banks_5_io_reads_2_en = 1'b1;
      end
    end
    if(when_BankedScratchMemory_l203_5) begin
      if(when_BankedScratchMemory_l206_45) begin
        banks_5_io_reads_2_en = 1'b1;
      end
    end
    if(when_BankedScratchMemory_l203_6) begin
      if(when_BankedScratchMemory_l206_53) begin
        banks_5_io_reads_2_en = 1'b1;
      end
    end
    if(when_BankedScratchMemory_l203_7) begin
      if(when_BankedScratchMemory_l206_61) begin
        banks_5_io_reads_2_en = 1'b1;
      end
    end
    if(when_BankedScratchMemory_l203_8) begin
      if(when_BankedScratchMemory_l206_69) begin
        banks_5_io_reads_2_en = 1'b1;
      end
    end
  end

  always @(*) begin
    banks_6_io_reads_0_addr = 8'h0;
    if(when_BankedScratchMemory_l160_6) begin
      banks_6_io_reads_0_addr = _zz_io_reads_0_addr;
    end
    if(when_BankedScratchMemory_l160_14) begin
      banks_6_io_reads_0_addr = _zz_io_reads_0_addr_1;
    end
    if(when_BankedScratchMemory_l160_22) begin
      banks_6_io_reads_0_addr = _zz_io_reads_0_addr_2;
    end
    if(when_BankedScratchMemory_l160_30) begin
      banks_6_io_reads_0_addr = _zz_io_reads_0_addr_3;
    end
    if(when_BankedScratchMemory_l160_38) begin
      banks_6_io_reads_0_addr = _zz_io_reads_0_addr_4;
    end
    if(when_BankedScratchMemory_l160_46) begin
      banks_6_io_reads_0_addr = _zz_io_reads_0_addr_5;
    end
    if(when_BankedScratchMemory_l160_54) begin
      banks_6_io_reads_0_addr = _zz_io_reads_0_addr_6;
    end
    if(when_BankedScratchMemory_l160_62) begin
      banks_6_io_reads_0_addr = _zz_io_reads_0_addr_7;
    end
  end

  always @(*) begin
    banks_6_io_reads_0_en = 1'b0;
    if(when_BankedScratchMemory_l160_6) begin
      banks_6_io_reads_0_en = io_valuReadEn_0_0;
    end
    if(when_BankedScratchMemory_l160_14) begin
      banks_6_io_reads_0_en = io_valuReadEn_0_1;
    end
    if(when_BankedScratchMemory_l160_22) begin
      banks_6_io_reads_0_en = io_valuReadEn_0_2;
    end
    if(when_BankedScratchMemory_l160_30) begin
      banks_6_io_reads_0_en = io_valuReadEn_0_3;
    end
    if(when_BankedScratchMemory_l160_38) begin
      banks_6_io_reads_0_en = io_valuReadEn_0_4;
    end
    if(when_BankedScratchMemory_l160_46) begin
      banks_6_io_reads_0_en = io_valuReadEn_0_5;
    end
    if(when_BankedScratchMemory_l160_54) begin
      banks_6_io_reads_0_en = io_valuReadEn_0_6;
    end
    if(when_BankedScratchMemory_l160_62) begin
      banks_6_io_reads_0_en = io_valuReadEn_0_7;
    end
  end

  always @(*) begin
    banks_6_io_reads_1_addr = 8'h0;
    if(when_BankedScratchMemory_l160_70) begin
      banks_6_io_reads_1_addr = _zz_io_reads_1_addr;
    end
    if(when_BankedScratchMemory_l160_78) begin
      banks_6_io_reads_1_addr = _zz_io_reads_1_addr_1;
    end
    if(when_BankedScratchMemory_l160_86) begin
      banks_6_io_reads_1_addr = _zz_io_reads_1_addr_2;
    end
    if(when_BankedScratchMemory_l160_94) begin
      banks_6_io_reads_1_addr = _zz_io_reads_1_addr_3;
    end
    if(when_BankedScratchMemory_l160_102) begin
      banks_6_io_reads_1_addr = _zz_io_reads_1_addr_4;
    end
    if(when_BankedScratchMemory_l160_110) begin
      banks_6_io_reads_1_addr = _zz_io_reads_1_addr_5;
    end
    if(when_BankedScratchMemory_l160_118) begin
      banks_6_io_reads_1_addr = _zz_io_reads_1_addr_6;
    end
    if(when_BankedScratchMemory_l160_126) begin
      banks_6_io_reads_1_addr = _zz_io_reads_1_addr_7;
    end
  end

  always @(*) begin
    banks_6_io_reads_1_en = 1'b0;
    if(when_BankedScratchMemory_l160_70) begin
      banks_6_io_reads_1_en = io_valuReadEn_1_0;
    end
    if(when_BankedScratchMemory_l160_78) begin
      banks_6_io_reads_1_en = io_valuReadEn_1_1;
    end
    if(when_BankedScratchMemory_l160_86) begin
      banks_6_io_reads_1_en = io_valuReadEn_1_2;
    end
    if(when_BankedScratchMemory_l160_94) begin
      banks_6_io_reads_1_en = io_valuReadEn_1_3;
    end
    if(when_BankedScratchMemory_l160_102) begin
      banks_6_io_reads_1_en = io_valuReadEn_1_4;
    end
    if(when_BankedScratchMemory_l160_110) begin
      banks_6_io_reads_1_en = io_valuReadEn_1_5;
    end
    if(when_BankedScratchMemory_l160_118) begin
      banks_6_io_reads_1_en = io_valuReadEn_1_6;
    end
    if(when_BankedScratchMemory_l160_126) begin
      banks_6_io_reads_1_en = io_valuReadEn_1_7;
    end
  end

  always @(*) begin
    banks_6_io_reads_2_addr = 8'h0;
    if(when_BankedScratchMemory_l203) begin
      if(when_BankedScratchMemory_l206_6) begin
        banks_6_io_reads_2_addr = scalarBankRow_0;
      end
    end
    if(when_BankedScratchMemory_l203_1) begin
      if(when_BankedScratchMemory_l206_14) begin
        banks_6_io_reads_2_addr = scalarBankRow_1;
      end
    end
    if(when_BankedScratchMemory_l203_2) begin
      if(when_BankedScratchMemory_l206_22) begin
        banks_6_io_reads_2_addr = scalarBankRow_2;
      end
    end
    if(when_BankedScratchMemory_l203_3) begin
      if(when_BankedScratchMemory_l206_30) begin
        banks_6_io_reads_2_addr = scalarBankRow_3;
      end
    end
    if(when_BankedScratchMemory_l203_4) begin
      if(when_BankedScratchMemory_l206_38) begin
        banks_6_io_reads_2_addr = scalarBankRow_4;
      end
    end
    if(when_BankedScratchMemory_l203_5) begin
      if(when_BankedScratchMemory_l206_46) begin
        banks_6_io_reads_2_addr = scalarBankRow_5;
      end
    end
    if(when_BankedScratchMemory_l203_6) begin
      if(when_BankedScratchMemory_l206_54) begin
        banks_6_io_reads_2_addr = scalarBankRow_6;
      end
    end
    if(when_BankedScratchMemory_l203_7) begin
      if(when_BankedScratchMemory_l206_62) begin
        banks_6_io_reads_2_addr = scalarBankRow_7;
      end
    end
    if(when_BankedScratchMemory_l203_8) begin
      if(when_BankedScratchMemory_l206_70) begin
        banks_6_io_reads_2_addr = scalarBankRow_8;
      end
    end
  end

  always @(*) begin
    banks_6_io_reads_2_en = 1'b0;
    if(when_BankedScratchMemory_l203) begin
      if(when_BankedScratchMemory_l206_6) begin
        banks_6_io_reads_2_en = 1'b1;
      end
    end
    if(when_BankedScratchMemory_l203_1) begin
      if(when_BankedScratchMemory_l206_14) begin
        banks_6_io_reads_2_en = 1'b1;
      end
    end
    if(when_BankedScratchMemory_l203_2) begin
      if(when_BankedScratchMemory_l206_22) begin
        banks_6_io_reads_2_en = 1'b1;
      end
    end
    if(when_BankedScratchMemory_l203_3) begin
      if(when_BankedScratchMemory_l206_30) begin
        banks_6_io_reads_2_en = 1'b1;
      end
    end
    if(when_BankedScratchMemory_l203_4) begin
      if(when_BankedScratchMemory_l206_38) begin
        banks_6_io_reads_2_en = 1'b1;
      end
    end
    if(when_BankedScratchMemory_l203_5) begin
      if(when_BankedScratchMemory_l206_46) begin
        banks_6_io_reads_2_en = 1'b1;
      end
    end
    if(when_BankedScratchMemory_l203_6) begin
      if(when_BankedScratchMemory_l206_54) begin
        banks_6_io_reads_2_en = 1'b1;
      end
    end
    if(when_BankedScratchMemory_l203_7) begin
      if(when_BankedScratchMemory_l206_62) begin
        banks_6_io_reads_2_en = 1'b1;
      end
    end
    if(when_BankedScratchMemory_l203_8) begin
      if(when_BankedScratchMemory_l206_70) begin
        banks_6_io_reads_2_en = 1'b1;
      end
    end
  end

  always @(*) begin
    banks_7_io_reads_0_addr = 8'h0;
    if(when_BankedScratchMemory_l160_7) begin
      banks_7_io_reads_0_addr = _zz_io_reads_0_addr;
    end
    if(when_BankedScratchMemory_l160_15) begin
      banks_7_io_reads_0_addr = _zz_io_reads_0_addr_1;
    end
    if(when_BankedScratchMemory_l160_23) begin
      banks_7_io_reads_0_addr = _zz_io_reads_0_addr_2;
    end
    if(when_BankedScratchMemory_l160_31) begin
      banks_7_io_reads_0_addr = _zz_io_reads_0_addr_3;
    end
    if(when_BankedScratchMemory_l160_39) begin
      banks_7_io_reads_0_addr = _zz_io_reads_0_addr_4;
    end
    if(when_BankedScratchMemory_l160_47) begin
      banks_7_io_reads_0_addr = _zz_io_reads_0_addr_5;
    end
    if(when_BankedScratchMemory_l160_55) begin
      banks_7_io_reads_0_addr = _zz_io_reads_0_addr_6;
    end
    if(when_BankedScratchMemory_l160_63) begin
      banks_7_io_reads_0_addr = _zz_io_reads_0_addr_7;
    end
  end

  always @(*) begin
    banks_7_io_reads_0_en = 1'b0;
    if(when_BankedScratchMemory_l160_7) begin
      banks_7_io_reads_0_en = io_valuReadEn_0_0;
    end
    if(when_BankedScratchMemory_l160_15) begin
      banks_7_io_reads_0_en = io_valuReadEn_0_1;
    end
    if(when_BankedScratchMemory_l160_23) begin
      banks_7_io_reads_0_en = io_valuReadEn_0_2;
    end
    if(when_BankedScratchMemory_l160_31) begin
      banks_7_io_reads_0_en = io_valuReadEn_0_3;
    end
    if(when_BankedScratchMemory_l160_39) begin
      banks_7_io_reads_0_en = io_valuReadEn_0_4;
    end
    if(when_BankedScratchMemory_l160_47) begin
      banks_7_io_reads_0_en = io_valuReadEn_0_5;
    end
    if(when_BankedScratchMemory_l160_55) begin
      banks_7_io_reads_0_en = io_valuReadEn_0_6;
    end
    if(when_BankedScratchMemory_l160_63) begin
      banks_7_io_reads_0_en = io_valuReadEn_0_7;
    end
  end

  always @(*) begin
    banks_7_io_reads_1_addr = 8'h0;
    if(when_BankedScratchMemory_l160_71) begin
      banks_7_io_reads_1_addr = _zz_io_reads_1_addr;
    end
    if(when_BankedScratchMemory_l160_79) begin
      banks_7_io_reads_1_addr = _zz_io_reads_1_addr_1;
    end
    if(when_BankedScratchMemory_l160_87) begin
      banks_7_io_reads_1_addr = _zz_io_reads_1_addr_2;
    end
    if(when_BankedScratchMemory_l160_95) begin
      banks_7_io_reads_1_addr = _zz_io_reads_1_addr_3;
    end
    if(when_BankedScratchMemory_l160_103) begin
      banks_7_io_reads_1_addr = _zz_io_reads_1_addr_4;
    end
    if(when_BankedScratchMemory_l160_111) begin
      banks_7_io_reads_1_addr = _zz_io_reads_1_addr_5;
    end
    if(when_BankedScratchMemory_l160_119) begin
      banks_7_io_reads_1_addr = _zz_io_reads_1_addr_6;
    end
    if(when_BankedScratchMemory_l160_127) begin
      banks_7_io_reads_1_addr = _zz_io_reads_1_addr_7;
    end
  end

  always @(*) begin
    banks_7_io_reads_1_en = 1'b0;
    if(when_BankedScratchMemory_l160_71) begin
      banks_7_io_reads_1_en = io_valuReadEn_1_0;
    end
    if(when_BankedScratchMemory_l160_79) begin
      banks_7_io_reads_1_en = io_valuReadEn_1_1;
    end
    if(when_BankedScratchMemory_l160_87) begin
      banks_7_io_reads_1_en = io_valuReadEn_1_2;
    end
    if(when_BankedScratchMemory_l160_95) begin
      banks_7_io_reads_1_en = io_valuReadEn_1_3;
    end
    if(when_BankedScratchMemory_l160_103) begin
      banks_7_io_reads_1_en = io_valuReadEn_1_4;
    end
    if(when_BankedScratchMemory_l160_111) begin
      banks_7_io_reads_1_en = io_valuReadEn_1_5;
    end
    if(when_BankedScratchMemory_l160_119) begin
      banks_7_io_reads_1_en = io_valuReadEn_1_6;
    end
    if(when_BankedScratchMemory_l160_127) begin
      banks_7_io_reads_1_en = io_valuReadEn_1_7;
    end
  end

  always @(*) begin
    banks_7_io_reads_2_addr = 8'h0;
    if(when_BankedScratchMemory_l203) begin
      if(when_BankedScratchMemory_l206_7) begin
        banks_7_io_reads_2_addr = scalarBankRow_0;
      end
    end
    if(when_BankedScratchMemory_l203_1) begin
      if(when_BankedScratchMemory_l206_15) begin
        banks_7_io_reads_2_addr = scalarBankRow_1;
      end
    end
    if(when_BankedScratchMemory_l203_2) begin
      if(when_BankedScratchMemory_l206_23) begin
        banks_7_io_reads_2_addr = scalarBankRow_2;
      end
    end
    if(when_BankedScratchMemory_l203_3) begin
      if(when_BankedScratchMemory_l206_31) begin
        banks_7_io_reads_2_addr = scalarBankRow_3;
      end
    end
    if(when_BankedScratchMemory_l203_4) begin
      if(when_BankedScratchMemory_l206_39) begin
        banks_7_io_reads_2_addr = scalarBankRow_4;
      end
    end
    if(when_BankedScratchMemory_l203_5) begin
      if(when_BankedScratchMemory_l206_47) begin
        banks_7_io_reads_2_addr = scalarBankRow_5;
      end
    end
    if(when_BankedScratchMemory_l203_6) begin
      if(when_BankedScratchMemory_l206_55) begin
        banks_7_io_reads_2_addr = scalarBankRow_6;
      end
    end
    if(when_BankedScratchMemory_l203_7) begin
      if(when_BankedScratchMemory_l206_63) begin
        banks_7_io_reads_2_addr = scalarBankRow_7;
      end
    end
    if(when_BankedScratchMemory_l203_8) begin
      if(when_BankedScratchMemory_l206_71) begin
        banks_7_io_reads_2_addr = scalarBankRow_8;
      end
    end
  end

  always @(*) begin
    banks_7_io_reads_2_en = 1'b0;
    if(when_BankedScratchMemory_l203) begin
      if(when_BankedScratchMemory_l206_7) begin
        banks_7_io_reads_2_en = 1'b1;
      end
    end
    if(when_BankedScratchMemory_l203_1) begin
      if(when_BankedScratchMemory_l206_15) begin
        banks_7_io_reads_2_en = 1'b1;
      end
    end
    if(when_BankedScratchMemory_l203_2) begin
      if(when_BankedScratchMemory_l206_23) begin
        banks_7_io_reads_2_en = 1'b1;
      end
    end
    if(when_BankedScratchMemory_l203_3) begin
      if(when_BankedScratchMemory_l206_31) begin
        banks_7_io_reads_2_en = 1'b1;
      end
    end
    if(when_BankedScratchMemory_l203_4) begin
      if(when_BankedScratchMemory_l206_39) begin
        banks_7_io_reads_2_en = 1'b1;
      end
    end
    if(when_BankedScratchMemory_l203_5) begin
      if(when_BankedScratchMemory_l206_47) begin
        banks_7_io_reads_2_en = 1'b1;
      end
    end
    if(when_BankedScratchMemory_l203_6) begin
      if(when_BankedScratchMemory_l206_55) begin
        banks_7_io_reads_2_en = 1'b1;
      end
    end
    if(when_BankedScratchMemory_l203_7) begin
      if(when_BankedScratchMemory_l206_63) begin
        banks_7_io_reads_2_en = 1'b1;
      end
    end
    if(when_BankedScratchMemory_l203_8) begin
      if(when_BankedScratchMemory_l206_71) begin
        banks_7_io_reads_2_en = 1'b1;
      end
    end
  end

  assign _zz_when_BankedScratchMemory_l160 = io_valuReadAddr_0_0[2 : 0];
  assign _zz_io_reads_0_addr = io_valuReadAddr_0_0[10 : 3];
  always @(*) begin
    _zz_io_valuReadData_0_0 = 32'h0;
    if(when_BankedScratchMemory_l160) begin
      _zz_io_valuReadData_0_0 = banks_0_io_reads_0_data;
    end
    if(when_BankedScratchMemory_l160_1) begin
      _zz_io_valuReadData_0_0 = banks_1_io_reads_0_data;
    end
    if(when_BankedScratchMemory_l160_2) begin
      _zz_io_valuReadData_0_0 = banks_2_io_reads_0_data;
    end
    if(when_BankedScratchMemory_l160_3) begin
      _zz_io_valuReadData_0_0 = banks_3_io_reads_0_data;
    end
    if(when_BankedScratchMemory_l160_4) begin
      _zz_io_valuReadData_0_0 = banks_4_io_reads_0_data;
    end
    if(when_BankedScratchMemory_l160_5) begin
      _zz_io_valuReadData_0_0 = banks_5_io_reads_0_data;
    end
    if(when_BankedScratchMemory_l160_6) begin
      _zz_io_valuReadData_0_0 = banks_6_io_reads_0_data;
    end
    if(when_BankedScratchMemory_l160_7) begin
      _zz_io_valuReadData_0_0 = banks_7_io_reads_0_data;
    end
  end

  assign when_BankedScratchMemory_l160 = (_zz_when_BankedScratchMemory_l160 == 3'b000);
  assign when_BankedScratchMemory_l160_1 = (_zz_when_BankedScratchMemory_l160 == 3'b001);
  assign when_BankedScratchMemory_l160_2 = (_zz_when_BankedScratchMemory_l160 == 3'b010);
  assign when_BankedScratchMemory_l160_3 = (_zz_when_BankedScratchMemory_l160 == 3'b011);
  assign when_BankedScratchMemory_l160_4 = (_zz_when_BankedScratchMemory_l160 == 3'b100);
  assign when_BankedScratchMemory_l160_5 = (_zz_when_BankedScratchMemory_l160 == 3'b101);
  assign when_BankedScratchMemory_l160_6 = (_zz_when_BankedScratchMemory_l160 == 3'b110);
  assign when_BankedScratchMemory_l160_7 = (_zz_when_BankedScratchMemory_l160 == 3'b111);
  assign io_valuReadData_0_0 = _zz_io_valuReadData_0_0;
  assign _zz_when_BankedScratchMemory_l160_1 = io_valuReadAddr_0_1[2 : 0];
  assign _zz_io_reads_0_addr_1 = io_valuReadAddr_0_1[10 : 3];
  always @(*) begin
    _zz_io_valuReadData_0_1 = 32'h0;
    if(when_BankedScratchMemory_l160_8) begin
      _zz_io_valuReadData_0_1 = banks_0_io_reads_0_data;
    end
    if(when_BankedScratchMemory_l160_9) begin
      _zz_io_valuReadData_0_1 = banks_1_io_reads_0_data;
    end
    if(when_BankedScratchMemory_l160_10) begin
      _zz_io_valuReadData_0_1 = banks_2_io_reads_0_data;
    end
    if(when_BankedScratchMemory_l160_11) begin
      _zz_io_valuReadData_0_1 = banks_3_io_reads_0_data;
    end
    if(when_BankedScratchMemory_l160_12) begin
      _zz_io_valuReadData_0_1 = banks_4_io_reads_0_data;
    end
    if(when_BankedScratchMemory_l160_13) begin
      _zz_io_valuReadData_0_1 = banks_5_io_reads_0_data;
    end
    if(when_BankedScratchMemory_l160_14) begin
      _zz_io_valuReadData_0_1 = banks_6_io_reads_0_data;
    end
    if(when_BankedScratchMemory_l160_15) begin
      _zz_io_valuReadData_0_1 = banks_7_io_reads_0_data;
    end
  end

  assign when_BankedScratchMemory_l160_8 = (_zz_when_BankedScratchMemory_l160_1 == 3'b000);
  assign when_BankedScratchMemory_l160_9 = (_zz_when_BankedScratchMemory_l160_1 == 3'b001);
  assign when_BankedScratchMemory_l160_10 = (_zz_when_BankedScratchMemory_l160_1 == 3'b010);
  assign when_BankedScratchMemory_l160_11 = (_zz_when_BankedScratchMemory_l160_1 == 3'b011);
  assign when_BankedScratchMemory_l160_12 = (_zz_when_BankedScratchMemory_l160_1 == 3'b100);
  assign when_BankedScratchMemory_l160_13 = (_zz_when_BankedScratchMemory_l160_1 == 3'b101);
  assign when_BankedScratchMemory_l160_14 = (_zz_when_BankedScratchMemory_l160_1 == 3'b110);
  assign when_BankedScratchMemory_l160_15 = (_zz_when_BankedScratchMemory_l160_1 == 3'b111);
  assign io_valuReadData_0_1 = _zz_io_valuReadData_0_1;
  assign _zz_when_BankedScratchMemory_l160_2 = io_valuReadAddr_0_2[2 : 0];
  assign _zz_io_reads_0_addr_2 = io_valuReadAddr_0_2[10 : 3];
  always @(*) begin
    _zz_io_valuReadData_0_2 = 32'h0;
    if(when_BankedScratchMemory_l160_16) begin
      _zz_io_valuReadData_0_2 = banks_0_io_reads_0_data;
    end
    if(when_BankedScratchMemory_l160_17) begin
      _zz_io_valuReadData_0_2 = banks_1_io_reads_0_data;
    end
    if(when_BankedScratchMemory_l160_18) begin
      _zz_io_valuReadData_0_2 = banks_2_io_reads_0_data;
    end
    if(when_BankedScratchMemory_l160_19) begin
      _zz_io_valuReadData_0_2 = banks_3_io_reads_0_data;
    end
    if(when_BankedScratchMemory_l160_20) begin
      _zz_io_valuReadData_0_2 = banks_4_io_reads_0_data;
    end
    if(when_BankedScratchMemory_l160_21) begin
      _zz_io_valuReadData_0_2 = banks_5_io_reads_0_data;
    end
    if(when_BankedScratchMemory_l160_22) begin
      _zz_io_valuReadData_0_2 = banks_6_io_reads_0_data;
    end
    if(when_BankedScratchMemory_l160_23) begin
      _zz_io_valuReadData_0_2 = banks_7_io_reads_0_data;
    end
  end

  assign when_BankedScratchMemory_l160_16 = (_zz_when_BankedScratchMemory_l160_2 == 3'b000);
  assign when_BankedScratchMemory_l160_17 = (_zz_when_BankedScratchMemory_l160_2 == 3'b001);
  assign when_BankedScratchMemory_l160_18 = (_zz_when_BankedScratchMemory_l160_2 == 3'b010);
  assign when_BankedScratchMemory_l160_19 = (_zz_when_BankedScratchMemory_l160_2 == 3'b011);
  assign when_BankedScratchMemory_l160_20 = (_zz_when_BankedScratchMemory_l160_2 == 3'b100);
  assign when_BankedScratchMemory_l160_21 = (_zz_when_BankedScratchMemory_l160_2 == 3'b101);
  assign when_BankedScratchMemory_l160_22 = (_zz_when_BankedScratchMemory_l160_2 == 3'b110);
  assign when_BankedScratchMemory_l160_23 = (_zz_when_BankedScratchMemory_l160_2 == 3'b111);
  assign io_valuReadData_0_2 = _zz_io_valuReadData_0_2;
  assign _zz_when_BankedScratchMemory_l160_3 = io_valuReadAddr_0_3[2 : 0];
  assign _zz_io_reads_0_addr_3 = io_valuReadAddr_0_3[10 : 3];
  always @(*) begin
    _zz_io_valuReadData_0_3 = 32'h0;
    if(when_BankedScratchMemory_l160_24) begin
      _zz_io_valuReadData_0_3 = banks_0_io_reads_0_data;
    end
    if(when_BankedScratchMemory_l160_25) begin
      _zz_io_valuReadData_0_3 = banks_1_io_reads_0_data;
    end
    if(when_BankedScratchMemory_l160_26) begin
      _zz_io_valuReadData_0_3 = banks_2_io_reads_0_data;
    end
    if(when_BankedScratchMemory_l160_27) begin
      _zz_io_valuReadData_0_3 = banks_3_io_reads_0_data;
    end
    if(when_BankedScratchMemory_l160_28) begin
      _zz_io_valuReadData_0_3 = banks_4_io_reads_0_data;
    end
    if(when_BankedScratchMemory_l160_29) begin
      _zz_io_valuReadData_0_3 = banks_5_io_reads_0_data;
    end
    if(when_BankedScratchMemory_l160_30) begin
      _zz_io_valuReadData_0_3 = banks_6_io_reads_0_data;
    end
    if(when_BankedScratchMemory_l160_31) begin
      _zz_io_valuReadData_0_3 = banks_7_io_reads_0_data;
    end
  end

  assign when_BankedScratchMemory_l160_24 = (_zz_when_BankedScratchMemory_l160_3 == 3'b000);
  assign when_BankedScratchMemory_l160_25 = (_zz_when_BankedScratchMemory_l160_3 == 3'b001);
  assign when_BankedScratchMemory_l160_26 = (_zz_when_BankedScratchMemory_l160_3 == 3'b010);
  assign when_BankedScratchMemory_l160_27 = (_zz_when_BankedScratchMemory_l160_3 == 3'b011);
  assign when_BankedScratchMemory_l160_28 = (_zz_when_BankedScratchMemory_l160_3 == 3'b100);
  assign when_BankedScratchMemory_l160_29 = (_zz_when_BankedScratchMemory_l160_3 == 3'b101);
  assign when_BankedScratchMemory_l160_30 = (_zz_when_BankedScratchMemory_l160_3 == 3'b110);
  assign when_BankedScratchMemory_l160_31 = (_zz_when_BankedScratchMemory_l160_3 == 3'b111);
  assign io_valuReadData_0_3 = _zz_io_valuReadData_0_3;
  assign _zz_when_BankedScratchMemory_l160_4 = io_valuReadAddr_0_4[2 : 0];
  assign _zz_io_reads_0_addr_4 = io_valuReadAddr_0_4[10 : 3];
  always @(*) begin
    _zz_io_valuReadData_0_4 = 32'h0;
    if(when_BankedScratchMemory_l160_32) begin
      _zz_io_valuReadData_0_4 = banks_0_io_reads_0_data;
    end
    if(when_BankedScratchMemory_l160_33) begin
      _zz_io_valuReadData_0_4 = banks_1_io_reads_0_data;
    end
    if(when_BankedScratchMemory_l160_34) begin
      _zz_io_valuReadData_0_4 = banks_2_io_reads_0_data;
    end
    if(when_BankedScratchMemory_l160_35) begin
      _zz_io_valuReadData_0_4 = banks_3_io_reads_0_data;
    end
    if(when_BankedScratchMemory_l160_36) begin
      _zz_io_valuReadData_0_4 = banks_4_io_reads_0_data;
    end
    if(when_BankedScratchMemory_l160_37) begin
      _zz_io_valuReadData_0_4 = banks_5_io_reads_0_data;
    end
    if(when_BankedScratchMemory_l160_38) begin
      _zz_io_valuReadData_0_4 = banks_6_io_reads_0_data;
    end
    if(when_BankedScratchMemory_l160_39) begin
      _zz_io_valuReadData_0_4 = banks_7_io_reads_0_data;
    end
  end

  assign when_BankedScratchMemory_l160_32 = (_zz_when_BankedScratchMemory_l160_4 == 3'b000);
  assign when_BankedScratchMemory_l160_33 = (_zz_when_BankedScratchMemory_l160_4 == 3'b001);
  assign when_BankedScratchMemory_l160_34 = (_zz_when_BankedScratchMemory_l160_4 == 3'b010);
  assign when_BankedScratchMemory_l160_35 = (_zz_when_BankedScratchMemory_l160_4 == 3'b011);
  assign when_BankedScratchMemory_l160_36 = (_zz_when_BankedScratchMemory_l160_4 == 3'b100);
  assign when_BankedScratchMemory_l160_37 = (_zz_when_BankedScratchMemory_l160_4 == 3'b101);
  assign when_BankedScratchMemory_l160_38 = (_zz_when_BankedScratchMemory_l160_4 == 3'b110);
  assign when_BankedScratchMemory_l160_39 = (_zz_when_BankedScratchMemory_l160_4 == 3'b111);
  assign io_valuReadData_0_4 = _zz_io_valuReadData_0_4;
  assign _zz_when_BankedScratchMemory_l160_5 = io_valuReadAddr_0_5[2 : 0];
  assign _zz_io_reads_0_addr_5 = io_valuReadAddr_0_5[10 : 3];
  always @(*) begin
    _zz_io_valuReadData_0_5 = 32'h0;
    if(when_BankedScratchMemory_l160_40) begin
      _zz_io_valuReadData_0_5 = banks_0_io_reads_0_data;
    end
    if(when_BankedScratchMemory_l160_41) begin
      _zz_io_valuReadData_0_5 = banks_1_io_reads_0_data;
    end
    if(when_BankedScratchMemory_l160_42) begin
      _zz_io_valuReadData_0_5 = banks_2_io_reads_0_data;
    end
    if(when_BankedScratchMemory_l160_43) begin
      _zz_io_valuReadData_0_5 = banks_3_io_reads_0_data;
    end
    if(when_BankedScratchMemory_l160_44) begin
      _zz_io_valuReadData_0_5 = banks_4_io_reads_0_data;
    end
    if(when_BankedScratchMemory_l160_45) begin
      _zz_io_valuReadData_0_5 = banks_5_io_reads_0_data;
    end
    if(when_BankedScratchMemory_l160_46) begin
      _zz_io_valuReadData_0_5 = banks_6_io_reads_0_data;
    end
    if(when_BankedScratchMemory_l160_47) begin
      _zz_io_valuReadData_0_5 = banks_7_io_reads_0_data;
    end
  end

  assign when_BankedScratchMemory_l160_40 = (_zz_when_BankedScratchMemory_l160_5 == 3'b000);
  assign when_BankedScratchMemory_l160_41 = (_zz_when_BankedScratchMemory_l160_5 == 3'b001);
  assign when_BankedScratchMemory_l160_42 = (_zz_when_BankedScratchMemory_l160_5 == 3'b010);
  assign when_BankedScratchMemory_l160_43 = (_zz_when_BankedScratchMemory_l160_5 == 3'b011);
  assign when_BankedScratchMemory_l160_44 = (_zz_when_BankedScratchMemory_l160_5 == 3'b100);
  assign when_BankedScratchMemory_l160_45 = (_zz_when_BankedScratchMemory_l160_5 == 3'b101);
  assign when_BankedScratchMemory_l160_46 = (_zz_when_BankedScratchMemory_l160_5 == 3'b110);
  assign when_BankedScratchMemory_l160_47 = (_zz_when_BankedScratchMemory_l160_5 == 3'b111);
  assign io_valuReadData_0_5 = _zz_io_valuReadData_0_5;
  assign _zz_when_BankedScratchMemory_l160_6 = io_valuReadAddr_0_6[2 : 0];
  assign _zz_io_reads_0_addr_6 = io_valuReadAddr_0_6[10 : 3];
  always @(*) begin
    _zz_io_valuReadData_0_6 = 32'h0;
    if(when_BankedScratchMemory_l160_48) begin
      _zz_io_valuReadData_0_6 = banks_0_io_reads_0_data;
    end
    if(when_BankedScratchMemory_l160_49) begin
      _zz_io_valuReadData_0_6 = banks_1_io_reads_0_data;
    end
    if(when_BankedScratchMemory_l160_50) begin
      _zz_io_valuReadData_0_6 = banks_2_io_reads_0_data;
    end
    if(when_BankedScratchMemory_l160_51) begin
      _zz_io_valuReadData_0_6 = banks_3_io_reads_0_data;
    end
    if(when_BankedScratchMemory_l160_52) begin
      _zz_io_valuReadData_0_6 = banks_4_io_reads_0_data;
    end
    if(when_BankedScratchMemory_l160_53) begin
      _zz_io_valuReadData_0_6 = banks_5_io_reads_0_data;
    end
    if(when_BankedScratchMemory_l160_54) begin
      _zz_io_valuReadData_0_6 = banks_6_io_reads_0_data;
    end
    if(when_BankedScratchMemory_l160_55) begin
      _zz_io_valuReadData_0_6 = banks_7_io_reads_0_data;
    end
  end

  assign when_BankedScratchMemory_l160_48 = (_zz_when_BankedScratchMemory_l160_6 == 3'b000);
  assign when_BankedScratchMemory_l160_49 = (_zz_when_BankedScratchMemory_l160_6 == 3'b001);
  assign when_BankedScratchMemory_l160_50 = (_zz_when_BankedScratchMemory_l160_6 == 3'b010);
  assign when_BankedScratchMemory_l160_51 = (_zz_when_BankedScratchMemory_l160_6 == 3'b011);
  assign when_BankedScratchMemory_l160_52 = (_zz_when_BankedScratchMemory_l160_6 == 3'b100);
  assign when_BankedScratchMemory_l160_53 = (_zz_when_BankedScratchMemory_l160_6 == 3'b101);
  assign when_BankedScratchMemory_l160_54 = (_zz_when_BankedScratchMemory_l160_6 == 3'b110);
  assign when_BankedScratchMemory_l160_55 = (_zz_when_BankedScratchMemory_l160_6 == 3'b111);
  assign io_valuReadData_0_6 = _zz_io_valuReadData_0_6;
  assign _zz_when_BankedScratchMemory_l160_7 = io_valuReadAddr_0_7[2 : 0];
  assign _zz_io_reads_0_addr_7 = io_valuReadAddr_0_7[10 : 3];
  always @(*) begin
    _zz_io_valuReadData_0_7 = 32'h0;
    if(when_BankedScratchMemory_l160_56) begin
      _zz_io_valuReadData_0_7 = banks_0_io_reads_0_data;
    end
    if(when_BankedScratchMemory_l160_57) begin
      _zz_io_valuReadData_0_7 = banks_1_io_reads_0_data;
    end
    if(when_BankedScratchMemory_l160_58) begin
      _zz_io_valuReadData_0_7 = banks_2_io_reads_0_data;
    end
    if(when_BankedScratchMemory_l160_59) begin
      _zz_io_valuReadData_0_7 = banks_3_io_reads_0_data;
    end
    if(when_BankedScratchMemory_l160_60) begin
      _zz_io_valuReadData_0_7 = banks_4_io_reads_0_data;
    end
    if(when_BankedScratchMemory_l160_61) begin
      _zz_io_valuReadData_0_7 = banks_5_io_reads_0_data;
    end
    if(when_BankedScratchMemory_l160_62) begin
      _zz_io_valuReadData_0_7 = banks_6_io_reads_0_data;
    end
    if(when_BankedScratchMemory_l160_63) begin
      _zz_io_valuReadData_0_7 = banks_7_io_reads_0_data;
    end
  end

  assign when_BankedScratchMemory_l160_56 = (_zz_when_BankedScratchMemory_l160_7 == 3'b000);
  assign when_BankedScratchMemory_l160_57 = (_zz_when_BankedScratchMemory_l160_7 == 3'b001);
  assign when_BankedScratchMemory_l160_58 = (_zz_when_BankedScratchMemory_l160_7 == 3'b010);
  assign when_BankedScratchMemory_l160_59 = (_zz_when_BankedScratchMemory_l160_7 == 3'b011);
  assign when_BankedScratchMemory_l160_60 = (_zz_when_BankedScratchMemory_l160_7 == 3'b100);
  assign when_BankedScratchMemory_l160_61 = (_zz_when_BankedScratchMemory_l160_7 == 3'b101);
  assign when_BankedScratchMemory_l160_62 = (_zz_when_BankedScratchMemory_l160_7 == 3'b110);
  assign when_BankedScratchMemory_l160_63 = (_zz_when_BankedScratchMemory_l160_7 == 3'b111);
  assign io_valuReadData_0_7 = _zz_io_valuReadData_0_7;
  assign _zz_when_BankedScratchMemory_l160_8 = io_valuReadAddr_1_0[2 : 0];
  assign _zz_io_reads_1_addr = io_valuReadAddr_1_0[10 : 3];
  always @(*) begin
    _zz_io_valuReadData_1_0 = 32'h0;
    if(when_BankedScratchMemory_l160_64) begin
      _zz_io_valuReadData_1_0 = banks_0_io_reads_1_data;
    end
    if(when_BankedScratchMemory_l160_65) begin
      _zz_io_valuReadData_1_0 = banks_1_io_reads_1_data;
    end
    if(when_BankedScratchMemory_l160_66) begin
      _zz_io_valuReadData_1_0 = banks_2_io_reads_1_data;
    end
    if(when_BankedScratchMemory_l160_67) begin
      _zz_io_valuReadData_1_0 = banks_3_io_reads_1_data;
    end
    if(when_BankedScratchMemory_l160_68) begin
      _zz_io_valuReadData_1_0 = banks_4_io_reads_1_data;
    end
    if(when_BankedScratchMemory_l160_69) begin
      _zz_io_valuReadData_1_0 = banks_5_io_reads_1_data;
    end
    if(when_BankedScratchMemory_l160_70) begin
      _zz_io_valuReadData_1_0 = banks_6_io_reads_1_data;
    end
    if(when_BankedScratchMemory_l160_71) begin
      _zz_io_valuReadData_1_0 = banks_7_io_reads_1_data;
    end
  end

  assign when_BankedScratchMemory_l160_64 = (_zz_when_BankedScratchMemory_l160_8 == 3'b000);
  assign when_BankedScratchMemory_l160_65 = (_zz_when_BankedScratchMemory_l160_8 == 3'b001);
  assign when_BankedScratchMemory_l160_66 = (_zz_when_BankedScratchMemory_l160_8 == 3'b010);
  assign when_BankedScratchMemory_l160_67 = (_zz_when_BankedScratchMemory_l160_8 == 3'b011);
  assign when_BankedScratchMemory_l160_68 = (_zz_when_BankedScratchMemory_l160_8 == 3'b100);
  assign when_BankedScratchMemory_l160_69 = (_zz_when_BankedScratchMemory_l160_8 == 3'b101);
  assign when_BankedScratchMemory_l160_70 = (_zz_when_BankedScratchMemory_l160_8 == 3'b110);
  assign when_BankedScratchMemory_l160_71 = (_zz_when_BankedScratchMemory_l160_8 == 3'b111);
  assign io_valuReadData_1_0 = _zz_io_valuReadData_1_0;
  assign _zz_when_BankedScratchMemory_l160_9 = io_valuReadAddr_1_1[2 : 0];
  assign _zz_io_reads_1_addr_1 = io_valuReadAddr_1_1[10 : 3];
  always @(*) begin
    _zz_io_valuReadData_1_1 = 32'h0;
    if(when_BankedScratchMemory_l160_72) begin
      _zz_io_valuReadData_1_1 = banks_0_io_reads_1_data;
    end
    if(when_BankedScratchMemory_l160_73) begin
      _zz_io_valuReadData_1_1 = banks_1_io_reads_1_data;
    end
    if(when_BankedScratchMemory_l160_74) begin
      _zz_io_valuReadData_1_1 = banks_2_io_reads_1_data;
    end
    if(when_BankedScratchMemory_l160_75) begin
      _zz_io_valuReadData_1_1 = banks_3_io_reads_1_data;
    end
    if(when_BankedScratchMemory_l160_76) begin
      _zz_io_valuReadData_1_1 = banks_4_io_reads_1_data;
    end
    if(when_BankedScratchMemory_l160_77) begin
      _zz_io_valuReadData_1_1 = banks_5_io_reads_1_data;
    end
    if(when_BankedScratchMemory_l160_78) begin
      _zz_io_valuReadData_1_1 = banks_6_io_reads_1_data;
    end
    if(when_BankedScratchMemory_l160_79) begin
      _zz_io_valuReadData_1_1 = banks_7_io_reads_1_data;
    end
  end

  assign when_BankedScratchMemory_l160_72 = (_zz_when_BankedScratchMemory_l160_9 == 3'b000);
  assign when_BankedScratchMemory_l160_73 = (_zz_when_BankedScratchMemory_l160_9 == 3'b001);
  assign when_BankedScratchMemory_l160_74 = (_zz_when_BankedScratchMemory_l160_9 == 3'b010);
  assign when_BankedScratchMemory_l160_75 = (_zz_when_BankedScratchMemory_l160_9 == 3'b011);
  assign when_BankedScratchMemory_l160_76 = (_zz_when_BankedScratchMemory_l160_9 == 3'b100);
  assign when_BankedScratchMemory_l160_77 = (_zz_when_BankedScratchMemory_l160_9 == 3'b101);
  assign when_BankedScratchMemory_l160_78 = (_zz_when_BankedScratchMemory_l160_9 == 3'b110);
  assign when_BankedScratchMemory_l160_79 = (_zz_when_BankedScratchMemory_l160_9 == 3'b111);
  assign io_valuReadData_1_1 = _zz_io_valuReadData_1_1;
  assign _zz_when_BankedScratchMemory_l160_10 = io_valuReadAddr_1_2[2 : 0];
  assign _zz_io_reads_1_addr_2 = io_valuReadAddr_1_2[10 : 3];
  always @(*) begin
    _zz_io_valuReadData_1_2 = 32'h0;
    if(when_BankedScratchMemory_l160_80) begin
      _zz_io_valuReadData_1_2 = banks_0_io_reads_1_data;
    end
    if(when_BankedScratchMemory_l160_81) begin
      _zz_io_valuReadData_1_2 = banks_1_io_reads_1_data;
    end
    if(when_BankedScratchMemory_l160_82) begin
      _zz_io_valuReadData_1_2 = banks_2_io_reads_1_data;
    end
    if(when_BankedScratchMemory_l160_83) begin
      _zz_io_valuReadData_1_2 = banks_3_io_reads_1_data;
    end
    if(when_BankedScratchMemory_l160_84) begin
      _zz_io_valuReadData_1_2 = banks_4_io_reads_1_data;
    end
    if(when_BankedScratchMemory_l160_85) begin
      _zz_io_valuReadData_1_2 = banks_5_io_reads_1_data;
    end
    if(when_BankedScratchMemory_l160_86) begin
      _zz_io_valuReadData_1_2 = banks_6_io_reads_1_data;
    end
    if(when_BankedScratchMemory_l160_87) begin
      _zz_io_valuReadData_1_2 = banks_7_io_reads_1_data;
    end
  end

  assign when_BankedScratchMemory_l160_80 = (_zz_when_BankedScratchMemory_l160_10 == 3'b000);
  assign when_BankedScratchMemory_l160_81 = (_zz_when_BankedScratchMemory_l160_10 == 3'b001);
  assign when_BankedScratchMemory_l160_82 = (_zz_when_BankedScratchMemory_l160_10 == 3'b010);
  assign when_BankedScratchMemory_l160_83 = (_zz_when_BankedScratchMemory_l160_10 == 3'b011);
  assign when_BankedScratchMemory_l160_84 = (_zz_when_BankedScratchMemory_l160_10 == 3'b100);
  assign when_BankedScratchMemory_l160_85 = (_zz_when_BankedScratchMemory_l160_10 == 3'b101);
  assign when_BankedScratchMemory_l160_86 = (_zz_when_BankedScratchMemory_l160_10 == 3'b110);
  assign when_BankedScratchMemory_l160_87 = (_zz_when_BankedScratchMemory_l160_10 == 3'b111);
  assign io_valuReadData_1_2 = _zz_io_valuReadData_1_2;
  assign _zz_when_BankedScratchMemory_l160_11 = io_valuReadAddr_1_3[2 : 0];
  assign _zz_io_reads_1_addr_3 = io_valuReadAddr_1_3[10 : 3];
  always @(*) begin
    _zz_io_valuReadData_1_3 = 32'h0;
    if(when_BankedScratchMemory_l160_88) begin
      _zz_io_valuReadData_1_3 = banks_0_io_reads_1_data;
    end
    if(when_BankedScratchMemory_l160_89) begin
      _zz_io_valuReadData_1_3 = banks_1_io_reads_1_data;
    end
    if(when_BankedScratchMemory_l160_90) begin
      _zz_io_valuReadData_1_3 = banks_2_io_reads_1_data;
    end
    if(when_BankedScratchMemory_l160_91) begin
      _zz_io_valuReadData_1_3 = banks_3_io_reads_1_data;
    end
    if(when_BankedScratchMemory_l160_92) begin
      _zz_io_valuReadData_1_3 = banks_4_io_reads_1_data;
    end
    if(when_BankedScratchMemory_l160_93) begin
      _zz_io_valuReadData_1_3 = banks_5_io_reads_1_data;
    end
    if(when_BankedScratchMemory_l160_94) begin
      _zz_io_valuReadData_1_3 = banks_6_io_reads_1_data;
    end
    if(when_BankedScratchMemory_l160_95) begin
      _zz_io_valuReadData_1_3 = banks_7_io_reads_1_data;
    end
  end

  assign when_BankedScratchMemory_l160_88 = (_zz_when_BankedScratchMemory_l160_11 == 3'b000);
  assign when_BankedScratchMemory_l160_89 = (_zz_when_BankedScratchMemory_l160_11 == 3'b001);
  assign when_BankedScratchMemory_l160_90 = (_zz_when_BankedScratchMemory_l160_11 == 3'b010);
  assign when_BankedScratchMemory_l160_91 = (_zz_when_BankedScratchMemory_l160_11 == 3'b011);
  assign when_BankedScratchMemory_l160_92 = (_zz_when_BankedScratchMemory_l160_11 == 3'b100);
  assign when_BankedScratchMemory_l160_93 = (_zz_when_BankedScratchMemory_l160_11 == 3'b101);
  assign when_BankedScratchMemory_l160_94 = (_zz_when_BankedScratchMemory_l160_11 == 3'b110);
  assign when_BankedScratchMemory_l160_95 = (_zz_when_BankedScratchMemory_l160_11 == 3'b111);
  assign io_valuReadData_1_3 = _zz_io_valuReadData_1_3;
  assign _zz_when_BankedScratchMemory_l160_12 = io_valuReadAddr_1_4[2 : 0];
  assign _zz_io_reads_1_addr_4 = io_valuReadAddr_1_4[10 : 3];
  always @(*) begin
    _zz_io_valuReadData_1_4 = 32'h0;
    if(when_BankedScratchMemory_l160_96) begin
      _zz_io_valuReadData_1_4 = banks_0_io_reads_1_data;
    end
    if(when_BankedScratchMemory_l160_97) begin
      _zz_io_valuReadData_1_4 = banks_1_io_reads_1_data;
    end
    if(when_BankedScratchMemory_l160_98) begin
      _zz_io_valuReadData_1_4 = banks_2_io_reads_1_data;
    end
    if(when_BankedScratchMemory_l160_99) begin
      _zz_io_valuReadData_1_4 = banks_3_io_reads_1_data;
    end
    if(when_BankedScratchMemory_l160_100) begin
      _zz_io_valuReadData_1_4 = banks_4_io_reads_1_data;
    end
    if(when_BankedScratchMemory_l160_101) begin
      _zz_io_valuReadData_1_4 = banks_5_io_reads_1_data;
    end
    if(when_BankedScratchMemory_l160_102) begin
      _zz_io_valuReadData_1_4 = banks_6_io_reads_1_data;
    end
    if(when_BankedScratchMemory_l160_103) begin
      _zz_io_valuReadData_1_4 = banks_7_io_reads_1_data;
    end
  end

  assign when_BankedScratchMemory_l160_96 = (_zz_when_BankedScratchMemory_l160_12 == 3'b000);
  assign when_BankedScratchMemory_l160_97 = (_zz_when_BankedScratchMemory_l160_12 == 3'b001);
  assign when_BankedScratchMemory_l160_98 = (_zz_when_BankedScratchMemory_l160_12 == 3'b010);
  assign when_BankedScratchMemory_l160_99 = (_zz_when_BankedScratchMemory_l160_12 == 3'b011);
  assign when_BankedScratchMemory_l160_100 = (_zz_when_BankedScratchMemory_l160_12 == 3'b100);
  assign when_BankedScratchMemory_l160_101 = (_zz_when_BankedScratchMemory_l160_12 == 3'b101);
  assign when_BankedScratchMemory_l160_102 = (_zz_when_BankedScratchMemory_l160_12 == 3'b110);
  assign when_BankedScratchMemory_l160_103 = (_zz_when_BankedScratchMemory_l160_12 == 3'b111);
  assign io_valuReadData_1_4 = _zz_io_valuReadData_1_4;
  assign _zz_when_BankedScratchMemory_l160_13 = io_valuReadAddr_1_5[2 : 0];
  assign _zz_io_reads_1_addr_5 = io_valuReadAddr_1_5[10 : 3];
  always @(*) begin
    _zz_io_valuReadData_1_5 = 32'h0;
    if(when_BankedScratchMemory_l160_104) begin
      _zz_io_valuReadData_1_5 = banks_0_io_reads_1_data;
    end
    if(when_BankedScratchMemory_l160_105) begin
      _zz_io_valuReadData_1_5 = banks_1_io_reads_1_data;
    end
    if(when_BankedScratchMemory_l160_106) begin
      _zz_io_valuReadData_1_5 = banks_2_io_reads_1_data;
    end
    if(when_BankedScratchMemory_l160_107) begin
      _zz_io_valuReadData_1_5 = banks_3_io_reads_1_data;
    end
    if(when_BankedScratchMemory_l160_108) begin
      _zz_io_valuReadData_1_5 = banks_4_io_reads_1_data;
    end
    if(when_BankedScratchMemory_l160_109) begin
      _zz_io_valuReadData_1_5 = banks_5_io_reads_1_data;
    end
    if(when_BankedScratchMemory_l160_110) begin
      _zz_io_valuReadData_1_5 = banks_6_io_reads_1_data;
    end
    if(when_BankedScratchMemory_l160_111) begin
      _zz_io_valuReadData_1_5 = banks_7_io_reads_1_data;
    end
  end

  assign when_BankedScratchMemory_l160_104 = (_zz_when_BankedScratchMemory_l160_13 == 3'b000);
  assign when_BankedScratchMemory_l160_105 = (_zz_when_BankedScratchMemory_l160_13 == 3'b001);
  assign when_BankedScratchMemory_l160_106 = (_zz_when_BankedScratchMemory_l160_13 == 3'b010);
  assign when_BankedScratchMemory_l160_107 = (_zz_when_BankedScratchMemory_l160_13 == 3'b011);
  assign when_BankedScratchMemory_l160_108 = (_zz_when_BankedScratchMemory_l160_13 == 3'b100);
  assign when_BankedScratchMemory_l160_109 = (_zz_when_BankedScratchMemory_l160_13 == 3'b101);
  assign when_BankedScratchMemory_l160_110 = (_zz_when_BankedScratchMemory_l160_13 == 3'b110);
  assign when_BankedScratchMemory_l160_111 = (_zz_when_BankedScratchMemory_l160_13 == 3'b111);
  assign io_valuReadData_1_5 = _zz_io_valuReadData_1_5;
  assign _zz_when_BankedScratchMemory_l160_14 = io_valuReadAddr_1_6[2 : 0];
  assign _zz_io_reads_1_addr_6 = io_valuReadAddr_1_6[10 : 3];
  always @(*) begin
    _zz_io_valuReadData_1_6 = 32'h0;
    if(when_BankedScratchMemory_l160_112) begin
      _zz_io_valuReadData_1_6 = banks_0_io_reads_1_data;
    end
    if(when_BankedScratchMemory_l160_113) begin
      _zz_io_valuReadData_1_6 = banks_1_io_reads_1_data;
    end
    if(when_BankedScratchMemory_l160_114) begin
      _zz_io_valuReadData_1_6 = banks_2_io_reads_1_data;
    end
    if(when_BankedScratchMemory_l160_115) begin
      _zz_io_valuReadData_1_6 = banks_3_io_reads_1_data;
    end
    if(when_BankedScratchMemory_l160_116) begin
      _zz_io_valuReadData_1_6 = banks_4_io_reads_1_data;
    end
    if(when_BankedScratchMemory_l160_117) begin
      _zz_io_valuReadData_1_6 = banks_5_io_reads_1_data;
    end
    if(when_BankedScratchMemory_l160_118) begin
      _zz_io_valuReadData_1_6 = banks_6_io_reads_1_data;
    end
    if(when_BankedScratchMemory_l160_119) begin
      _zz_io_valuReadData_1_6 = banks_7_io_reads_1_data;
    end
  end

  assign when_BankedScratchMemory_l160_112 = (_zz_when_BankedScratchMemory_l160_14 == 3'b000);
  assign when_BankedScratchMemory_l160_113 = (_zz_when_BankedScratchMemory_l160_14 == 3'b001);
  assign when_BankedScratchMemory_l160_114 = (_zz_when_BankedScratchMemory_l160_14 == 3'b010);
  assign when_BankedScratchMemory_l160_115 = (_zz_when_BankedScratchMemory_l160_14 == 3'b011);
  assign when_BankedScratchMemory_l160_116 = (_zz_when_BankedScratchMemory_l160_14 == 3'b100);
  assign when_BankedScratchMemory_l160_117 = (_zz_when_BankedScratchMemory_l160_14 == 3'b101);
  assign when_BankedScratchMemory_l160_118 = (_zz_when_BankedScratchMemory_l160_14 == 3'b110);
  assign when_BankedScratchMemory_l160_119 = (_zz_when_BankedScratchMemory_l160_14 == 3'b111);
  assign io_valuReadData_1_6 = _zz_io_valuReadData_1_6;
  assign _zz_when_BankedScratchMemory_l160_15 = io_valuReadAddr_1_7[2 : 0];
  assign _zz_io_reads_1_addr_7 = io_valuReadAddr_1_7[10 : 3];
  always @(*) begin
    _zz_io_valuReadData_1_7 = 32'h0;
    if(when_BankedScratchMemory_l160_120) begin
      _zz_io_valuReadData_1_7 = banks_0_io_reads_1_data;
    end
    if(when_BankedScratchMemory_l160_121) begin
      _zz_io_valuReadData_1_7 = banks_1_io_reads_1_data;
    end
    if(when_BankedScratchMemory_l160_122) begin
      _zz_io_valuReadData_1_7 = banks_2_io_reads_1_data;
    end
    if(when_BankedScratchMemory_l160_123) begin
      _zz_io_valuReadData_1_7 = banks_3_io_reads_1_data;
    end
    if(when_BankedScratchMemory_l160_124) begin
      _zz_io_valuReadData_1_7 = banks_4_io_reads_1_data;
    end
    if(when_BankedScratchMemory_l160_125) begin
      _zz_io_valuReadData_1_7 = banks_5_io_reads_1_data;
    end
    if(when_BankedScratchMemory_l160_126) begin
      _zz_io_valuReadData_1_7 = banks_6_io_reads_1_data;
    end
    if(when_BankedScratchMemory_l160_127) begin
      _zz_io_valuReadData_1_7 = banks_7_io_reads_1_data;
    end
  end

  assign when_BankedScratchMemory_l160_120 = (_zz_when_BankedScratchMemory_l160_15 == 3'b000);
  assign when_BankedScratchMemory_l160_121 = (_zz_when_BankedScratchMemory_l160_15 == 3'b001);
  assign when_BankedScratchMemory_l160_122 = (_zz_when_BankedScratchMemory_l160_15 == 3'b010);
  assign when_BankedScratchMemory_l160_123 = (_zz_when_BankedScratchMemory_l160_15 == 3'b011);
  assign when_BankedScratchMemory_l160_124 = (_zz_when_BankedScratchMemory_l160_15 == 3'b100);
  assign when_BankedScratchMemory_l160_125 = (_zz_when_BankedScratchMemory_l160_15 == 3'b101);
  assign when_BankedScratchMemory_l160_126 = (_zz_when_BankedScratchMemory_l160_15 == 3'b110);
  assign when_BankedScratchMemory_l160_127 = (_zz_when_BankedScratchMemory_l160_15 == 3'b111);
  assign io_valuReadData_1_7 = _zz_io_valuReadData_1_7;
  always @(*) begin
    io_conflict = 1'b0;
    if(when_BankedScratchMemory_l213) begin
      io_conflict = 1'b1;
    end
    if(when_BankedScratchMemory_l213_1) begin
      io_conflict = 1'b1;
    end
    if(when_BankedScratchMemory_l213_2) begin
      io_conflict = 1'b1;
    end
    if(when_BankedScratchMemory_l213_3) begin
      io_conflict = 1'b1;
    end
    if(when_BankedScratchMemory_l213_4) begin
      io_conflict = 1'b1;
    end
    if(when_BankedScratchMemory_l213_5) begin
      io_conflict = 1'b1;
    end
    if(when_BankedScratchMemory_l213_6) begin
      io_conflict = 1'b1;
    end
    if(when_BankedScratchMemory_l213_7) begin
      io_conflict = 1'b1;
    end
    if(when_BankedScratchMemory_l213_8) begin
      io_conflict = 1'b1;
    end
  end

  assign scalarBankReq_0 = io_scalarReadAddr_0[2 : 0];
  assign scalarBankRow_0 = io_scalarReadAddr_0[10 : 3];
  always @(*) begin
    io_scalarReadData_0 = 32'h0;
    if(when_BankedScratchMemory_l222) begin
      io_scalarReadData_0 = banks_0_io_reads_2_data;
    end
    if(when_BankedScratchMemory_l222_1) begin
      io_scalarReadData_0 = banks_1_io_reads_2_data;
    end
    if(when_BankedScratchMemory_l222_2) begin
      io_scalarReadData_0 = banks_2_io_reads_2_data;
    end
    if(when_BankedScratchMemory_l222_3) begin
      io_scalarReadData_0 = banks_3_io_reads_2_data;
    end
    if(when_BankedScratchMemory_l222_4) begin
      io_scalarReadData_0 = banks_4_io_reads_2_data;
    end
    if(when_BankedScratchMemory_l222_5) begin
      io_scalarReadData_0 = banks_5_io_reads_2_data;
    end
    if(when_BankedScratchMemory_l222_6) begin
      io_scalarReadData_0 = banks_6_io_reads_2_data;
    end
    if(when_BankedScratchMemory_l222_7) begin
      io_scalarReadData_0 = banks_7_io_reads_2_data;
    end
  end

  assign scalarBankReq_1 = io_scalarReadAddr_1[2 : 0];
  assign scalarBankRow_1 = io_scalarReadAddr_1[10 : 3];
  always @(*) begin
    io_scalarReadData_1 = 32'h0;
    if(when_BankedScratchMemory_l222_8) begin
      io_scalarReadData_1 = banks_0_io_reads_2_data;
    end
    if(when_BankedScratchMemory_l222_9) begin
      io_scalarReadData_1 = banks_1_io_reads_2_data;
    end
    if(when_BankedScratchMemory_l222_10) begin
      io_scalarReadData_1 = banks_2_io_reads_2_data;
    end
    if(when_BankedScratchMemory_l222_11) begin
      io_scalarReadData_1 = banks_3_io_reads_2_data;
    end
    if(when_BankedScratchMemory_l222_12) begin
      io_scalarReadData_1 = banks_4_io_reads_2_data;
    end
    if(when_BankedScratchMemory_l222_13) begin
      io_scalarReadData_1 = banks_5_io_reads_2_data;
    end
    if(when_BankedScratchMemory_l222_14) begin
      io_scalarReadData_1 = banks_6_io_reads_2_data;
    end
    if(when_BankedScratchMemory_l222_15) begin
      io_scalarReadData_1 = banks_7_io_reads_2_data;
    end
  end

  assign scalarBankReq_2 = io_scalarReadAddr_2[2 : 0];
  assign scalarBankRow_2 = io_scalarReadAddr_2[10 : 3];
  always @(*) begin
    io_scalarReadData_2 = 32'h0;
    if(when_BankedScratchMemory_l222_16) begin
      io_scalarReadData_2 = banks_0_io_reads_2_data;
    end
    if(when_BankedScratchMemory_l222_17) begin
      io_scalarReadData_2 = banks_1_io_reads_2_data;
    end
    if(when_BankedScratchMemory_l222_18) begin
      io_scalarReadData_2 = banks_2_io_reads_2_data;
    end
    if(when_BankedScratchMemory_l222_19) begin
      io_scalarReadData_2 = banks_3_io_reads_2_data;
    end
    if(when_BankedScratchMemory_l222_20) begin
      io_scalarReadData_2 = banks_4_io_reads_2_data;
    end
    if(when_BankedScratchMemory_l222_21) begin
      io_scalarReadData_2 = banks_5_io_reads_2_data;
    end
    if(when_BankedScratchMemory_l222_22) begin
      io_scalarReadData_2 = banks_6_io_reads_2_data;
    end
    if(when_BankedScratchMemory_l222_23) begin
      io_scalarReadData_2 = banks_7_io_reads_2_data;
    end
  end

  assign scalarBankReq_3 = io_scalarReadAddr_3[2 : 0];
  assign scalarBankRow_3 = io_scalarReadAddr_3[10 : 3];
  always @(*) begin
    io_scalarReadData_3 = 32'h0;
    if(when_BankedScratchMemory_l222_24) begin
      io_scalarReadData_3 = banks_0_io_reads_2_data;
    end
    if(when_BankedScratchMemory_l222_25) begin
      io_scalarReadData_3 = banks_1_io_reads_2_data;
    end
    if(when_BankedScratchMemory_l222_26) begin
      io_scalarReadData_3 = banks_2_io_reads_2_data;
    end
    if(when_BankedScratchMemory_l222_27) begin
      io_scalarReadData_3 = banks_3_io_reads_2_data;
    end
    if(when_BankedScratchMemory_l222_28) begin
      io_scalarReadData_3 = banks_4_io_reads_2_data;
    end
    if(when_BankedScratchMemory_l222_29) begin
      io_scalarReadData_3 = banks_5_io_reads_2_data;
    end
    if(when_BankedScratchMemory_l222_30) begin
      io_scalarReadData_3 = banks_6_io_reads_2_data;
    end
    if(when_BankedScratchMemory_l222_31) begin
      io_scalarReadData_3 = banks_7_io_reads_2_data;
    end
  end

  assign scalarBankReq_4 = io_scalarReadAddr_4[2 : 0];
  assign scalarBankRow_4 = io_scalarReadAddr_4[10 : 3];
  always @(*) begin
    io_scalarReadData_4 = 32'h0;
    if(when_BankedScratchMemory_l222_32) begin
      io_scalarReadData_4 = banks_0_io_reads_2_data;
    end
    if(when_BankedScratchMemory_l222_33) begin
      io_scalarReadData_4 = banks_1_io_reads_2_data;
    end
    if(when_BankedScratchMemory_l222_34) begin
      io_scalarReadData_4 = banks_2_io_reads_2_data;
    end
    if(when_BankedScratchMemory_l222_35) begin
      io_scalarReadData_4 = banks_3_io_reads_2_data;
    end
    if(when_BankedScratchMemory_l222_36) begin
      io_scalarReadData_4 = banks_4_io_reads_2_data;
    end
    if(when_BankedScratchMemory_l222_37) begin
      io_scalarReadData_4 = banks_5_io_reads_2_data;
    end
    if(when_BankedScratchMemory_l222_38) begin
      io_scalarReadData_4 = banks_6_io_reads_2_data;
    end
    if(when_BankedScratchMemory_l222_39) begin
      io_scalarReadData_4 = banks_7_io_reads_2_data;
    end
  end

  assign scalarBankReq_5 = io_scalarReadAddr_5[2 : 0];
  assign scalarBankRow_5 = io_scalarReadAddr_5[10 : 3];
  always @(*) begin
    io_scalarReadData_5 = 32'h0;
    if(when_BankedScratchMemory_l222_40) begin
      io_scalarReadData_5 = banks_0_io_reads_2_data;
    end
    if(when_BankedScratchMemory_l222_41) begin
      io_scalarReadData_5 = banks_1_io_reads_2_data;
    end
    if(when_BankedScratchMemory_l222_42) begin
      io_scalarReadData_5 = banks_2_io_reads_2_data;
    end
    if(when_BankedScratchMemory_l222_43) begin
      io_scalarReadData_5 = banks_3_io_reads_2_data;
    end
    if(when_BankedScratchMemory_l222_44) begin
      io_scalarReadData_5 = banks_4_io_reads_2_data;
    end
    if(when_BankedScratchMemory_l222_45) begin
      io_scalarReadData_5 = banks_5_io_reads_2_data;
    end
    if(when_BankedScratchMemory_l222_46) begin
      io_scalarReadData_5 = banks_6_io_reads_2_data;
    end
    if(when_BankedScratchMemory_l222_47) begin
      io_scalarReadData_5 = banks_7_io_reads_2_data;
    end
  end

  assign scalarBankReq_6 = io_scalarReadAddr_6[2 : 0];
  assign scalarBankRow_6 = io_scalarReadAddr_6[10 : 3];
  always @(*) begin
    io_scalarReadData_6 = 32'h0;
    if(when_BankedScratchMemory_l222_48) begin
      io_scalarReadData_6 = banks_0_io_reads_2_data;
    end
    if(when_BankedScratchMemory_l222_49) begin
      io_scalarReadData_6 = banks_1_io_reads_2_data;
    end
    if(when_BankedScratchMemory_l222_50) begin
      io_scalarReadData_6 = banks_2_io_reads_2_data;
    end
    if(when_BankedScratchMemory_l222_51) begin
      io_scalarReadData_6 = banks_3_io_reads_2_data;
    end
    if(when_BankedScratchMemory_l222_52) begin
      io_scalarReadData_6 = banks_4_io_reads_2_data;
    end
    if(when_BankedScratchMemory_l222_53) begin
      io_scalarReadData_6 = banks_5_io_reads_2_data;
    end
    if(when_BankedScratchMemory_l222_54) begin
      io_scalarReadData_6 = banks_6_io_reads_2_data;
    end
    if(when_BankedScratchMemory_l222_55) begin
      io_scalarReadData_6 = banks_7_io_reads_2_data;
    end
  end

  assign scalarBankReq_7 = io_scalarReadAddr_7[2 : 0];
  assign scalarBankRow_7 = io_scalarReadAddr_7[10 : 3];
  always @(*) begin
    io_scalarReadData_7 = 32'h0;
    if(when_BankedScratchMemory_l222_56) begin
      io_scalarReadData_7 = banks_0_io_reads_2_data;
    end
    if(when_BankedScratchMemory_l222_57) begin
      io_scalarReadData_7 = banks_1_io_reads_2_data;
    end
    if(when_BankedScratchMemory_l222_58) begin
      io_scalarReadData_7 = banks_2_io_reads_2_data;
    end
    if(when_BankedScratchMemory_l222_59) begin
      io_scalarReadData_7 = banks_3_io_reads_2_data;
    end
    if(when_BankedScratchMemory_l222_60) begin
      io_scalarReadData_7 = banks_4_io_reads_2_data;
    end
    if(when_BankedScratchMemory_l222_61) begin
      io_scalarReadData_7 = banks_5_io_reads_2_data;
    end
    if(when_BankedScratchMemory_l222_62) begin
      io_scalarReadData_7 = banks_6_io_reads_2_data;
    end
    if(when_BankedScratchMemory_l222_63) begin
      io_scalarReadData_7 = banks_7_io_reads_2_data;
    end
  end

  assign scalarBankReq_8 = io_scalarReadAddr_8[2 : 0];
  assign scalarBankRow_8 = io_scalarReadAddr_8[10 : 3];
  always @(*) begin
    io_scalarReadData_8 = 32'h0;
    if(when_BankedScratchMemory_l222_64) begin
      io_scalarReadData_8 = banks_0_io_reads_2_data;
    end
    if(when_BankedScratchMemory_l222_65) begin
      io_scalarReadData_8 = banks_1_io_reads_2_data;
    end
    if(when_BankedScratchMemory_l222_66) begin
      io_scalarReadData_8 = banks_2_io_reads_2_data;
    end
    if(when_BankedScratchMemory_l222_67) begin
      io_scalarReadData_8 = banks_3_io_reads_2_data;
    end
    if(when_BankedScratchMemory_l222_68) begin
      io_scalarReadData_8 = banks_4_io_reads_2_data;
    end
    if(when_BankedScratchMemory_l222_69) begin
      io_scalarReadData_8 = banks_5_io_reads_2_data;
    end
    if(when_BankedScratchMemory_l222_70) begin
      io_scalarReadData_8 = banks_6_io_reads_2_data;
    end
    if(when_BankedScratchMemory_l222_71) begin
      io_scalarReadData_8 = banks_7_io_reads_2_data;
    end
  end

  assign _zz_when_BankedScratchMemory_l203 = 1'b0;
  assign when_BankedScratchMemory_l203 = (io_scalarReadEn_0 && (! _zz_when_BankedScratchMemory_l203));
  assign when_BankedScratchMemory_l206 = (scalarBankReq_0 == 3'b000);
  assign when_BankedScratchMemory_l206_1 = (scalarBankReq_0 == 3'b001);
  assign when_BankedScratchMemory_l206_2 = (scalarBankReq_0 == 3'b010);
  assign when_BankedScratchMemory_l206_3 = (scalarBankReq_0 == 3'b011);
  assign when_BankedScratchMemory_l206_4 = (scalarBankReq_0 == 3'b100);
  assign when_BankedScratchMemory_l206_5 = (scalarBankReq_0 == 3'b101);
  assign when_BankedScratchMemory_l206_6 = (scalarBankReq_0 == 3'b110);
  assign when_BankedScratchMemory_l206_7 = (scalarBankReq_0 == 3'b111);
  assign when_BankedScratchMemory_l213 = (io_scalarReadEn_0 && _zz_when_BankedScratchMemory_l203);
  assign _zz_when_BankedScratchMemory_l203_1 = (io_scalarReadEn_0 && (scalarBankReq_0 == scalarBankReq_1));
  assign when_BankedScratchMemory_l203_1 = (io_scalarReadEn_1 && (! _zz_when_BankedScratchMemory_l203_1));
  assign when_BankedScratchMemory_l206_8 = (scalarBankReq_1 == 3'b000);
  assign when_BankedScratchMemory_l206_9 = (scalarBankReq_1 == 3'b001);
  assign when_BankedScratchMemory_l206_10 = (scalarBankReq_1 == 3'b010);
  assign when_BankedScratchMemory_l206_11 = (scalarBankReq_1 == 3'b011);
  assign when_BankedScratchMemory_l206_12 = (scalarBankReq_1 == 3'b100);
  assign when_BankedScratchMemory_l206_13 = (scalarBankReq_1 == 3'b101);
  assign when_BankedScratchMemory_l206_14 = (scalarBankReq_1 == 3'b110);
  assign when_BankedScratchMemory_l206_15 = (scalarBankReq_1 == 3'b111);
  assign when_BankedScratchMemory_l213_1 = (io_scalarReadEn_1 && _zz_when_BankedScratchMemory_l203_1);
  assign _zz_when_BankedScratchMemory_l203_2 = ((io_scalarReadEn_0 && (scalarBankReq_0 == scalarBankReq_2)) || (io_scalarReadEn_1 && (scalarBankReq_1 == scalarBankReq_2)));
  assign when_BankedScratchMemory_l203_2 = (io_scalarReadEn_2 && (! _zz_when_BankedScratchMemory_l203_2));
  assign when_BankedScratchMemory_l206_16 = (scalarBankReq_2 == 3'b000);
  assign when_BankedScratchMemory_l206_17 = (scalarBankReq_2 == 3'b001);
  assign when_BankedScratchMemory_l206_18 = (scalarBankReq_2 == 3'b010);
  assign when_BankedScratchMemory_l206_19 = (scalarBankReq_2 == 3'b011);
  assign when_BankedScratchMemory_l206_20 = (scalarBankReq_2 == 3'b100);
  assign when_BankedScratchMemory_l206_21 = (scalarBankReq_2 == 3'b101);
  assign when_BankedScratchMemory_l206_22 = (scalarBankReq_2 == 3'b110);
  assign when_BankedScratchMemory_l206_23 = (scalarBankReq_2 == 3'b111);
  assign when_BankedScratchMemory_l213_2 = (io_scalarReadEn_2 && _zz_when_BankedScratchMemory_l203_2);
  assign _zz_when_BankedScratchMemory_l203_3 = (((io_scalarReadEn_0 && (scalarBankReq_0 == scalarBankReq_3)) || (io_scalarReadEn_1 && (scalarBankReq_1 == scalarBankReq_3))) || (io_scalarReadEn_2 && (scalarBankReq_2 == scalarBankReq_3)));
  assign when_BankedScratchMemory_l203_3 = (io_scalarReadEn_3 && (! _zz_when_BankedScratchMemory_l203_3));
  assign when_BankedScratchMemory_l206_24 = (scalarBankReq_3 == 3'b000);
  assign when_BankedScratchMemory_l206_25 = (scalarBankReq_3 == 3'b001);
  assign when_BankedScratchMemory_l206_26 = (scalarBankReq_3 == 3'b010);
  assign when_BankedScratchMemory_l206_27 = (scalarBankReq_3 == 3'b011);
  assign when_BankedScratchMemory_l206_28 = (scalarBankReq_3 == 3'b100);
  assign when_BankedScratchMemory_l206_29 = (scalarBankReq_3 == 3'b101);
  assign when_BankedScratchMemory_l206_30 = (scalarBankReq_3 == 3'b110);
  assign when_BankedScratchMemory_l206_31 = (scalarBankReq_3 == 3'b111);
  assign when_BankedScratchMemory_l213_3 = (io_scalarReadEn_3 && _zz_when_BankedScratchMemory_l203_3);
  assign _zz_when_BankedScratchMemory_l203_4 = ((((io_scalarReadEn_0 && (scalarBankReq_0 == scalarBankReq_4)) || (io_scalarReadEn_1 && (scalarBankReq_1 == scalarBankReq_4))) || (io_scalarReadEn_2 && (scalarBankReq_2 == scalarBankReq_4))) || (io_scalarReadEn_3 && (scalarBankReq_3 == scalarBankReq_4)));
  assign when_BankedScratchMemory_l203_4 = (io_scalarReadEn_4 && (! _zz_when_BankedScratchMemory_l203_4));
  assign when_BankedScratchMemory_l206_32 = (scalarBankReq_4 == 3'b000);
  assign when_BankedScratchMemory_l206_33 = (scalarBankReq_4 == 3'b001);
  assign when_BankedScratchMemory_l206_34 = (scalarBankReq_4 == 3'b010);
  assign when_BankedScratchMemory_l206_35 = (scalarBankReq_4 == 3'b011);
  assign when_BankedScratchMemory_l206_36 = (scalarBankReq_4 == 3'b100);
  assign when_BankedScratchMemory_l206_37 = (scalarBankReq_4 == 3'b101);
  assign when_BankedScratchMemory_l206_38 = (scalarBankReq_4 == 3'b110);
  assign when_BankedScratchMemory_l206_39 = (scalarBankReq_4 == 3'b111);
  assign when_BankedScratchMemory_l213_4 = (io_scalarReadEn_4 && _zz_when_BankedScratchMemory_l203_4);
  assign _zz_when_BankedScratchMemory_l203_5 = (((((io_scalarReadEn_0 && (scalarBankReq_0 == scalarBankReq_5)) || (io_scalarReadEn_1 && (scalarBankReq_1 == scalarBankReq_5))) || (io_scalarReadEn_2 && (scalarBankReq_2 == scalarBankReq_5))) || (io_scalarReadEn_3 && (scalarBankReq_3 == scalarBankReq_5))) || (io_scalarReadEn_4 && (scalarBankReq_4 == scalarBankReq_5)));
  assign when_BankedScratchMemory_l203_5 = (io_scalarReadEn_5 && (! _zz_when_BankedScratchMemory_l203_5));
  assign when_BankedScratchMemory_l206_40 = (scalarBankReq_5 == 3'b000);
  assign when_BankedScratchMemory_l206_41 = (scalarBankReq_5 == 3'b001);
  assign when_BankedScratchMemory_l206_42 = (scalarBankReq_5 == 3'b010);
  assign when_BankedScratchMemory_l206_43 = (scalarBankReq_5 == 3'b011);
  assign when_BankedScratchMemory_l206_44 = (scalarBankReq_5 == 3'b100);
  assign when_BankedScratchMemory_l206_45 = (scalarBankReq_5 == 3'b101);
  assign when_BankedScratchMemory_l206_46 = (scalarBankReq_5 == 3'b110);
  assign when_BankedScratchMemory_l206_47 = (scalarBankReq_5 == 3'b111);
  assign when_BankedScratchMemory_l213_5 = (io_scalarReadEn_5 && _zz_when_BankedScratchMemory_l203_5);
  assign _zz_when_BankedScratchMemory_l203_6 = ((((((io_scalarReadEn_0 && (scalarBankReq_0 == scalarBankReq_6)) || (io_scalarReadEn_1 && (scalarBankReq_1 == scalarBankReq_6))) || (io_scalarReadEn_2 && (scalarBankReq_2 == scalarBankReq_6))) || (io_scalarReadEn_3 && (scalarBankReq_3 == scalarBankReq_6))) || (io_scalarReadEn_4 && (scalarBankReq_4 == scalarBankReq_6))) || (io_scalarReadEn_5 && (scalarBankReq_5 == scalarBankReq_6)));
  assign when_BankedScratchMemory_l203_6 = (io_scalarReadEn_6 && (! _zz_when_BankedScratchMemory_l203_6));
  assign when_BankedScratchMemory_l206_48 = (scalarBankReq_6 == 3'b000);
  assign when_BankedScratchMemory_l206_49 = (scalarBankReq_6 == 3'b001);
  assign when_BankedScratchMemory_l206_50 = (scalarBankReq_6 == 3'b010);
  assign when_BankedScratchMemory_l206_51 = (scalarBankReq_6 == 3'b011);
  assign when_BankedScratchMemory_l206_52 = (scalarBankReq_6 == 3'b100);
  assign when_BankedScratchMemory_l206_53 = (scalarBankReq_6 == 3'b101);
  assign when_BankedScratchMemory_l206_54 = (scalarBankReq_6 == 3'b110);
  assign when_BankedScratchMemory_l206_55 = (scalarBankReq_6 == 3'b111);
  assign when_BankedScratchMemory_l213_6 = (io_scalarReadEn_6 && _zz_when_BankedScratchMemory_l203_6);
  assign _zz_when_BankedScratchMemory_l203_7 = (((((((io_scalarReadEn_0 && _zz__zz_when_BankedScratchMemory_l203_7) || (io_scalarReadEn_1 && _zz__zz_when_BankedScratchMemory_l203_7_1)) || (io_scalarReadEn_2 && (scalarBankReq_2 == scalarBankReq_7))) || (io_scalarReadEn_3 && (scalarBankReq_3 == scalarBankReq_7))) || (io_scalarReadEn_4 && (scalarBankReq_4 == scalarBankReq_7))) || (io_scalarReadEn_5 && (scalarBankReq_5 == scalarBankReq_7))) || (io_scalarReadEn_6 && (scalarBankReq_6 == scalarBankReq_7)));
  assign when_BankedScratchMemory_l203_7 = (io_scalarReadEn_7 && (! _zz_when_BankedScratchMemory_l203_7));
  assign when_BankedScratchMemory_l206_56 = (scalarBankReq_7 == 3'b000);
  assign when_BankedScratchMemory_l206_57 = (scalarBankReq_7 == 3'b001);
  assign when_BankedScratchMemory_l206_58 = (scalarBankReq_7 == 3'b010);
  assign when_BankedScratchMemory_l206_59 = (scalarBankReq_7 == 3'b011);
  assign when_BankedScratchMemory_l206_60 = (scalarBankReq_7 == 3'b100);
  assign when_BankedScratchMemory_l206_61 = (scalarBankReq_7 == 3'b101);
  assign when_BankedScratchMemory_l206_62 = (scalarBankReq_7 == 3'b110);
  assign when_BankedScratchMemory_l206_63 = (scalarBankReq_7 == 3'b111);
  assign when_BankedScratchMemory_l213_7 = (io_scalarReadEn_7 && _zz_when_BankedScratchMemory_l203_7);
  assign _zz_when_BankedScratchMemory_l203_8 = (((((((_zz__zz_when_BankedScratchMemory_l203_8 || _zz__zz_when_BankedScratchMemory_l203_8_1) || (io_scalarReadEn_2 && _zz__zz_when_BankedScratchMemory_l203_8_2)) || (io_scalarReadEn_3 && (scalarBankReq_3 == scalarBankReq_8))) || (io_scalarReadEn_4 && (scalarBankReq_4 == scalarBankReq_8))) || (io_scalarReadEn_5 && (scalarBankReq_5 == scalarBankReq_8))) || (io_scalarReadEn_6 && (scalarBankReq_6 == scalarBankReq_8))) || (io_scalarReadEn_7 && (scalarBankReq_7 == scalarBankReq_8)));
  assign when_BankedScratchMemory_l203_8 = (io_scalarReadEn_8 && (! _zz_when_BankedScratchMemory_l203_8));
  assign when_BankedScratchMemory_l206_64 = (scalarBankReq_8 == 3'b000);
  assign when_BankedScratchMemory_l206_65 = (scalarBankReq_8 == 3'b001);
  assign when_BankedScratchMemory_l206_66 = (scalarBankReq_8 == 3'b010);
  assign when_BankedScratchMemory_l206_67 = (scalarBankReq_8 == 3'b011);
  assign when_BankedScratchMemory_l206_68 = (scalarBankReq_8 == 3'b100);
  assign when_BankedScratchMemory_l206_69 = (scalarBankReq_8 == 3'b101);
  assign when_BankedScratchMemory_l206_70 = (scalarBankReq_8 == 3'b110);
  assign when_BankedScratchMemory_l206_71 = (scalarBankReq_8 == 3'b111);
  assign when_BankedScratchMemory_l213_8 = (io_scalarReadEn_8 && _zz_when_BankedScratchMemory_l203_8);
  assign when_BankedScratchMemory_l222 = (scalarBankReq_0 == 3'b000);
  assign when_BankedScratchMemory_l222_1 = (scalarBankReq_0 == 3'b001);
  assign when_BankedScratchMemory_l222_2 = (scalarBankReq_0 == 3'b010);
  assign when_BankedScratchMemory_l222_3 = (scalarBankReq_0 == 3'b011);
  assign when_BankedScratchMemory_l222_4 = (scalarBankReq_0 == 3'b100);
  assign when_BankedScratchMemory_l222_5 = (scalarBankReq_0 == 3'b101);
  assign when_BankedScratchMemory_l222_6 = (scalarBankReq_0 == 3'b110);
  assign when_BankedScratchMemory_l222_7 = (scalarBankReq_0 == 3'b111);
  assign when_BankedScratchMemory_l222_8 = (scalarBankReq_1 == 3'b000);
  assign when_BankedScratchMemory_l222_9 = (scalarBankReq_1 == 3'b001);
  assign when_BankedScratchMemory_l222_10 = (scalarBankReq_1 == 3'b010);
  assign when_BankedScratchMemory_l222_11 = (scalarBankReq_1 == 3'b011);
  assign when_BankedScratchMemory_l222_12 = (scalarBankReq_1 == 3'b100);
  assign when_BankedScratchMemory_l222_13 = (scalarBankReq_1 == 3'b101);
  assign when_BankedScratchMemory_l222_14 = (scalarBankReq_1 == 3'b110);
  assign when_BankedScratchMemory_l222_15 = (scalarBankReq_1 == 3'b111);
  assign when_BankedScratchMemory_l222_16 = (scalarBankReq_2 == 3'b000);
  assign when_BankedScratchMemory_l222_17 = (scalarBankReq_2 == 3'b001);
  assign when_BankedScratchMemory_l222_18 = (scalarBankReq_2 == 3'b010);
  assign when_BankedScratchMemory_l222_19 = (scalarBankReq_2 == 3'b011);
  assign when_BankedScratchMemory_l222_20 = (scalarBankReq_2 == 3'b100);
  assign when_BankedScratchMemory_l222_21 = (scalarBankReq_2 == 3'b101);
  assign when_BankedScratchMemory_l222_22 = (scalarBankReq_2 == 3'b110);
  assign when_BankedScratchMemory_l222_23 = (scalarBankReq_2 == 3'b111);
  assign when_BankedScratchMemory_l222_24 = (scalarBankReq_3 == 3'b000);
  assign when_BankedScratchMemory_l222_25 = (scalarBankReq_3 == 3'b001);
  assign when_BankedScratchMemory_l222_26 = (scalarBankReq_3 == 3'b010);
  assign when_BankedScratchMemory_l222_27 = (scalarBankReq_3 == 3'b011);
  assign when_BankedScratchMemory_l222_28 = (scalarBankReq_3 == 3'b100);
  assign when_BankedScratchMemory_l222_29 = (scalarBankReq_3 == 3'b101);
  assign when_BankedScratchMemory_l222_30 = (scalarBankReq_3 == 3'b110);
  assign when_BankedScratchMemory_l222_31 = (scalarBankReq_3 == 3'b111);
  assign when_BankedScratchMemory_l222_32 = (scalarBankReq_4 == 3'b000);
  assign when_BankedScratchMemory_l222_33 = (scalarBankReq_4 == 3'b001);
  assign when_BankedScratchMemory_l222_34 = (scalarBankReq_4 == 3'b010);
  assign when_BankedScratchMemory_l222_35 = (scalarBankReq_4 == 3'b011);
  assign when_BankedScratchMemory_l222_36 = (scalarBankReq_4 == 3'b100);
  assign when_BankedScratchMemory_l222_37 = (scalarBankReq_4 == 3'b101);
  assign when_BankedScratchMemory_l222_38 = (scalarBankReq_4 == 3'b110);
  assign when_BankedScratchMemory_l222_39 = (scalarBankReq_4 == 3'b111);
  assign when_BankedScratchMemory_l222_40 = (scalarBankReq_5 == 3'b000);
  assign when_BankedScratchMemory_l222_41 = (scalarBankReq_5 == 3'b001);
  assign when_BankedScratchMemory_l222_42 = (scalarBankReq_5 == 3'b010);
  assign when_BankedScratchMemory_l222_43 = (scalarBankReq_5 == 3'b011);
  assign when_BankedScratchMemory_l222_44 = (scalarBankReq_5 == 3'b100);
  assign when_BankedScratchMemory_l222_45 = (scalarBankReq_5 == 3'b101);
  assign when_BankedScratchMemory_l222_46 = (scalarBankReq_5 == 3'b110);
  assign when_BankedScratchMemory_l222_47 = (scalarBankReq_5 == 3'b111);
  assign when_BankedScratchMemory_l222_48 = (scalarBankReq_6 == 3'b000);
  assign when_BankedScratchMemory_l222_49 = (scalarBankReq_6 == 3'b001);
  assign when_BankedScratchMemory_l222_50 = (scalarBankReq_6 == 3'b010);
  assign when_BankedScratchMemory_l222_51 = (scalarBankReq_6 == 3'b011);
  assign when_BankedScratchMemory_l222_52 = (scalarBankReq_6 == 3'b100);
  assign when_BankedScratchMemory_l222_53 = (scalarBankReq_6 == 3'b101);
  assign when_BankedScratchMemory_l222_54 = (scalarBankReq_6 == 3'b110);
  assign when_BankedScratchMemory_l222_55 = (scalarBankReq_6 == 3'b111);
  assign when_BankedScratchMemory_l222_56 = (scalarBankReq_7 == 3'b000);
  assign when_BankedScratchMemory_l222_57 = (scalarBankReq_7 == 3'b001);
  assign when_BankedScratchMemory_l222_58 = (scalarBankReq_7 == 3'b010);
  assign when_BankedScratchMemory_l222_59 = (scalarBankReq_7 == 3'b011);
  assign when_BankedScratchMemory_l222_60 = (scalarBankReq_7 == 3'b100);
  assign when_BankedScratchMemory_l222_61 = (scalarBankReq_7 == 3'b101);
  assign when_BankedScratchMemory_l222_62 = (scalarBankReq_7 == 3'b110);
  assign when_BankedScratchMemory_l222_63 = (scalarBankReq_7 == 3'b111);
  assign when_BankedScratchMemory_l222_64 = (scalarBankReq_8 == 3'b000);
  assign when_BankedScratchMemory_l222_65 = (scalarBankReq_8 == 3'b001);
  assign when_BankedScratchMemory_l222_66 = (scalarBankReq_8 == 3'b010);
  assign when_BankedScratchMemory_l222_67 = (scalarBankReq_8 == 3'b011);
  assign when_BankedScratchMemory_l222_68 = (scalarBankReq_8 == 3'b100);
  assign when_BankedScratchMemory_l222_69 = (scalarBankReq_8 == 3'b101);
  assign when_BankedScratchMemory_l222_70 = (scalarBankReq_8 == 3'b110);
  assign when_BankedScratchMemory_l222_71 = (scalarBankReq_8 == 3'b111);
  always @(*) begin
    banks_0_io_write_en = 1'b0;
    if(io_writeEn_0) begin
      if(when_BankedScratchMemory_l242) begin
        banks_0_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_1) begin
      if(when_BankedScratchMemory_l242_8) begin
        banks_0_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_2) begin
      if(when_BankedScratchMemory_l242_16) begin
        banks_0_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_3) begin
      if(when_BankedScratchMemory_l242_24) begin
        banks_0_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_4) begin
      if(when_BankedScratchMemory_l242_32) begin
        banks_0_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_5) begin
      if(when_BankedScratchMemory_l242_40) begin
        banks_0_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_6) begin
      if(when_BankedScratchMemory_l242_48) begin
        banks_0_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_7) begin
      if(when_BankedScratchMemory_l242_56) begin
        banks_0_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_8) begin
      if(when_BankedScratchMemory_l242_64) begin
        banks_0_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_9) begin
      if(when_BankedScratchMemory_l242_72) begin
        banks_0_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_10) begin
      if(when_BankedScratchMemory_l242_80) begin
        banks_0_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_11) begin
      if(when_BankedScratchMemory_l242_88) begin
        banks_0_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_12) begin
      if(when_BankedScratchMemory_l242_96) begin
        banks_0_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_13) begin
      if(when_BankedScratchMemory_l242_104) begin
        banks_0_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_14) begin
      if(when_BankedScratchMemory_l242_112) begin
        banks_0_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_15) begin
      if(when_BankedScratchMemory_l242_120) begin
        banks_0_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_16) begin
      if(when_BankedScratchMemory_l242_128) begin
        banks_0_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_17) begin
      if(when_BankedScratchMemory_l242_136) begin
        banks_0_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_18) begin
      if(when_BankedScratchMemory_l242_144) begin
        banks_0_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_19) begin
      if(when_BankedScratchMemory_l242_152) begin
        banks_0_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_20) begin
      if(when_BankedScratchMemory_l242_160) begin
        banks_0_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_21) begin
      if(when_BankedScratchMemory_l242_168) begin
        banks_0_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_22) begin
      if(when_BankedScratchMemory_l242_176) begin
        banks_0_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_23) begin
      if(when_BankedScratchMemory_l242_184) begin
        banks_0_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_24) begin
      if(when_BankedScratchMemory_l242_192) begin
        banks_0_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_25) begin
      if(when_BankedScratchMemory_l242_200) begin
        banks_0_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_26) begin
      if(when_BankedScratchMemory_l242_208) begin
        banks_0_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_27) begin
      if(when_BankedScratchMemory_l242_216) begin
        banks_0_io_write_en = 1'b1;
      end
    end
  end

  always @(*) begin
    banks_0_io_write_addr = 8'h0;
    if(io_writeEn_0) begin
      if(when_BankedScratchMemory_l242) begin
        banks_0_io_write_addr = _zz_io_write_addr;
      end
    end
    if(io_writeEn_1) begin
      if(when_BankedScratchMemory_l242_8) begin
        banks_0_io_write_addr = _zz_io_write_addr_1;
      end
    end
    if(io_writeEn_2) begin
      if(when_BankedScratchMemory_l242_16) begin
        banks_0_io_write_addr = _zz_io_write_addr_2;
      end
    end
    if(io_writeEn_3) begin
      if(when_BankedScratchMemory_l242_24) begin
        banks_0_io_write_addr = _zz_io_write_addr_3;
      end
    end
    if(io_writeEn_4) begin
      if(when_BankedScratchMemory_l242_32) begin
        banks_0_io_write_addr = _zz_io_write_addr_4;
      end
    end
    if(io_writeEn_5) begin
      if(when_BankedScratchMemory_l242_40) begin
        banks_0_io_write_addr = _zz_io_write_addr_5;
      end
    end
    if(io_writeEn_6) begin
      if(when_BankedScratchMemory_l242_48) begin
        banks_0_io_write_addr = _zz_io_write_addr_6;
      end
    end
    if(io_writeEn_7) begin
      if(when_BankedScratchMemory_l242_56) begin
        banks_0_io_write_addr = _zz_io_write_addr_7;
      end
    end
    if(io_writeEn_8) begin
      if(when_BankedScratchMemory_l242_64) begin
        banks_0_io_write_addr = _zz_io_write_addr_8;
      end
    end
    if(io_writeEn_9) begin
      if(when_BankedScratchMemory_l242_72) begin
        banks_0_io_write_addr = _zz_io_write_addr_9;
      end
    end
    if(io_writeEn_10) begin
      if(when_BankedScratchMemory_l242_80) begin
        banks_0_io_write_addr = _zz_io_write_addr_10;
      end
    end
    if(io_writeEn_11) begin
      if(when_BankedScratchMemory_l242_88) begin
        banks_0_io_write_addr = _zz_io_write_addr_11;
      end
    end
    if(io_writeEn_12) begin
      if(when_BankedScratchMemory_l242_96) begin
        banks_0_io_write_addr = _zz_io_write_addr_12;
      end
    end
    if(io_writeEn_13) begin
      if(when_BankedScratchMemory_l242_104) begin
        banks_0_io_write_addr = _zz_io_write_addr_13;
      end
    end
    if(io_writeEn_14) begin
      if(when_BankedScratchMemory_l242_112) begin
        banks_0_io_write_addr = _zz_io_write_addr_14;
      end
    end
    if(io_writeEn_15) begin
      if(when_BankedScratchMemory_l242_120) begin
        banks_0_io_write_addr = _zz_io_write_addr_15;
      end
    end
    if(io_writeEn_16) begin
      if(when_BankedScratchMemory_l242_128) begin
        banks_0_io_write_addr = _zz_io_write_addr_16;
      end
    end
    if(io_writeEn_17) begin
      if(when_BankedScratchMemory_l242_136) begin
        banks_0_io_write_addr = _zz_io_write_addr_17;
      end
    end
    if(io_writeEn_18) begin
      if(when_BankedScratchMemory_l242_144) begin
        banks_0_io_write_addr = _zz_io_write_addr_18;
      end
    end
    if(io_writeEn_19) begin
      if(when_BankedScratchMemory_l242_152) begin
        banks_0_io_write_addr = _zz_io_write_addr_19;
      end
    end
    if(io_writeEn_20) begin
      if(when_BankedScratchMemory_l242_160) begin
        banks_0_io_write_addr = _zz_io_write_addr_20;
      end
    end
    if(io_writeEn_21) begin
      if(when_BankedScratchMemory_l242_168) begin
        banks_0_io_write_addr = _zz_io_write_addr_21;
      end
    end
    if(io_writeEn_22) begin
      if(when_BankedScratchMemory_l242_176) begin
        banks_0_io_write_addr = _zz_io_write_addr_22;
      end
    end
    if(io_writeEn_23) begin
      if(when_BankedScratchMemory_l242_184) begin
        banks_0_io_write_addr = _zz_io_write_addr_23;
      end
    end
    if(io_writeEn_24) begin
      if(when_BankedScratchMemory_l242_192) begin
        banks_0_io_write_addr = _zz_io_write_addr_24;
      end
    end
    if(io_writeEn_25) begin
      if(when_BankedScratchMemory_l242_200) begin
        banks_0_io_write_addr = _zz_io_write_addr_25;
      end
    end
    if(io_writeEn_26) begin
      if(when_BankedScratchMemory_l242_208) begin
        banks_0_io_write_addr = _zz_io_write_addr_26;
      end
    end
    if(io_writeEn_27) begin
      if(when_BankedScratchMemory_l242_216) begin
        banks_0_io_write_addr = _zz_io_write_addr_27;
      end
    end
  end

  always @(*) begin
    banks_0_io_write_data = 32'h0;
    if(io_writeEn_0) begin
      if(when_BankedScratchMemory_l242) begin
        banks_0_io_write_data = io_writeData_0;
      end
    end
    if(io_writeEn_1) begin
      if(when_BankedScratchMemory_l242_8) begin
        banks_0_io_write_data = io_writeData_1;
      end
    end
    if(io_writeEn_2) begin
      if(when_BankedScratchMemory_l242_16) begin
        banks_0_io_write_data = io_writeData_2;
      end
    end
    if(io_writeEn_3) begin
      if(when_BankedScratchMemory_l242_24) begin
        banks_0_io_write_data = io_writeData_3;
      end
    end
    if(io_writeEn_4) begin
      if(when_BankedScratchMemory_l242_32) begin
        banks_0_io_write_data = io_writeData_4;
      end
    end
    if(io_writeEn_5) begin
      if(when_BankedScratchMemory_l242_40) begin
        banks_0_io_write_data = io_writeData_5;
      end
    end
    if(io_writeEn_6) begin
      if(when_BankedScratchMemory_l242_48) begin
        banks_0_io_write_data = io_writeData_6;
      end
    end
    if(io_writeEn_7) begin
      if(when_BankedScratchMemory_l242_56) begin
        banks_0_io_write_data = io_writeData_7;
      end
    end
    if(io_writeEn_8) begin
      if(when_BankedScratchMemory_l242_64) begin
        banks_0_io_write_data = io_writeData_8;
      end
    end
    if(io_writeEn_9) begin
      if(when_BankedScratchMemory_l242_72) begin
        banks_0_io_write_data = io_writeData_9;
      end
    end
    if(io_writeEn_10) begin
      if(when_BankedScratchMemory_l242_80) begin
        banks_0_io_write_data = io_writeData_10;
      end
    end
    if(io_writeEn_11) begin
      if(when_BankedScratchMemory_l242_88) begin
        banks_0_io_write_data = io_writeData_11;
      end
    end
    if(io_writeEn_12) begin
      if(when_BankedScratchMemory_l242_96) begin
        banks_0_io_write_data = io_writeData_12;
      end
    end
    if(io_writeEn_13) begin
      if(when_BankedScratchMemory_l242_104) begin
        banks_0_io_write_data = io_writeData_13;
      end
    end
    if(io_writeEn_14) begin
      if(when_BankedScratchMemory_l242_112) begin
        banks_0_io_write_data = io_writeData_14;
      end
    end
    if(io_writeEn_15) begin
      if(when_BankedScratchMemory_l242_120) begin
        banks_0_io_write_data = io_writeData_15;
      end
    end
    if(io_writeEn_16) begin
      if(when_BankedScratchMemory_l242_128) begin
        banks_0_io_write_data = io_writeData_16;
      end
    end
    if(io_writeEn_17) begin
      if(when_BankedScratchMemory_l242_136) begin
        banks_0_io_write_data = io_writeData_17;
      end
    end
    if(io_writeEn_18) begin
      if(when_BankedScratchMemory_l242_144) begin
        banks_0_io_write_data = io_writeData_18;
      end
    end
    if(io_writeEn_19) begin
      if(when_BankedScratchMemory_l242_152) begin
        banks_0_io_write_data = io_writeData_19;
      end
    end
    if(io_writeEn_20) begin
      if(when_BankedScratchMemory_l242_160) begin
        banks_0_io_write_data = io_writeData_20;
      end
    end
    if(io_writeEn_21) begin
      if(when_BankedScratchMemory_l242_168) begin
        banks_0_io_write_data = io_writeData_21;
      end
    end
    if(io_writeEn_22) begin
      if(when_BankedScratchMemory_l242_176) begin
        banks_0_io_write_data = io_writeData_22;
      end
    end
    if(io_writeEn_23) begin
      if(when_BankedScratchMemory_l242_184) begin
        banks_0_io_write_data = io_writeData_23;
      end
    end
    if(io_writeEn_24) begin
      if(when_BankedScratchMemory_l242_192) begin
        banks_0_io_write_data = io_writeData_24;
      end
    end
    if(io_writeEn_25) begin
      if(when_BankedScratchMemory_l242_200) begin
        banks_0_io_write_data = io_writeData_25;
      end
    end
    if(io_writeEn_26) begin
      if(when_BankedScratchMemory_l242_208) begin
        banks_0_io_write_data = io_writeData_26;
      end
    end
    if(io_writeEn_27) begin
      if(when_BankedScratchMemory_l242_216) begin
        banks_0_io_write_data = io_writeData_27;
      end
    end
  end

  always @(*) begin
    banks_1_io_write_en = 1'b0;
    if(io_writeEn_0) begin
      if(when_BankedScratchMemory_l242_1) begin
        banks_1_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_1) begin
      if(when_BankedScratchMemory_l242_9) begin
        banks_1_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_2) begin
      if(when_BankedScratchMemory_l242_17) begin
        banks_1_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_3) begin
      if(when_BankedScratchMemory_l242_25) begin
        banks_1_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_4) begin
      if(when_BankedScratchMemory_l242_33) begin
        banks_1_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_5) begin
      if(when_BankedScratchMemory_l242_41) begin
        banks_1_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_6) begin
      if(when_BankedScratchMemory_l242_49) begin
        banks_1_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_7) begin
      if(when_BankedScratchMemory_l242_57) begin
        banks_1_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_8) begin
      if(when_BankedScratchMemory_l242_65) begin
        banks_1_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_9) begin
      if(when_BankedScratchMemory_l242_73) begin
        banks_1_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_10) begin
      if(when_BankedScratchMemory_l242_81) begin
        banks_1_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_11) begin
      if(when_BankedScratchMemory_l242_89) begin
        banks_1_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_12) begin
      if(when_BankedScratchMemory_l242_97) begin
        banks_1_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_13) begin
      if(when_BankedScratchMemory_l242_105) begin
        banks_1_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_14) begin
      if(when_BankedScratchMemory_l242_113) begin
        banks_1_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_15) begin
      if(when_BankedScratchMemory_l242_121) begin
        banks_1_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_16) begin
      if(when_BankedScratchMemory_l242_129) begin
        banks_1_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_17) begin
      if(when_BankedScratchMemory_l242_137) begin
        banks_1_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_18) begin
      if(when_BankedScratchMemory_l242_145) begin
        banks_1_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_19) begin
      if(when_BankedScratchMemory_l242_153) begin
        banks_1_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_20) begin
      if(when_BankedScratchMemory_l242_161) begin
        banks_1_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_21) begin
      if(when_BankedScratchMemory_l242_169) begin
        banks_1_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_22) begin
      if(when_BankedScratchMemory_l242_177) begin
        banks_1_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_23) begin
      if(when_BankedScratchMemory_l242_185) begin
        banks_1_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_24) begin
      if(when_BankedScratchMemory_l242_193) begin
        banks_1_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_25) begin
      if(when_BankedScratchMemory_l242_201) begin
        banks_1_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_26) begin
      if(when_BankedScratchMemory_l242_209) begin
        banks_1_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_27) begin
      if(when_BankedScratchMemory_l242_217) begin
        banks_1_io_write_en = 1'b1;
      end
    end
  end

  always @(*) begin
    banks_1_io_write_addr = 8'h0;
    if(io_writeEn_0) begin
      if(when_BankedScratchMemory_l242_1) begin
        banks_1_io_write_addr = _zz_io_write_addr;
      end
    end
    if(io_writeEn_1) begin
      if(when_BankedScratchMemory_l242_9) begin
        banks_1_io_write_addr = _zz_io_write_addr_1;
      end
    end
    if(io_writeEn_2) begin
      if(when_BankedScratchMemory_l242_17) begin
        banks_1_io_write_addr = _zz_io_write_addr_2;
      end
    end
    if(io_writeEn_3) begin
      if(when_BankedScratchMemory_l242_25) begin
        banks_1_io_write_addr = _zz_io_write_addr_3;
      end
    end
    if(io_writeEn_4) begin
      if(when_BankedScratchMemory_l242_33) begin
        banks_1_io_write_addr = _zz_io_write_addr_4;
      end
    end
    if(io_writeEn_5) begin
      if(when_BankedScratchMemory_l242_41) begin
        banks_1_io_write_addr = _zz_io_write_addr_5;
      end
    end
    if(io_writeEn_6) begin
      if(when_BankedScratchMemory_l242_49) begin
        banks_1_io_write_addr = _zz_io_write_addr_6;
      end
    end
    if(io_writeEn_7) begin
      if(when_BankedScratchMemory_l242_57) begin
        banks_1_io_write_addr = _zz_io_write_addr_7;
      end
    end
    if(io_writeEn_8) begin
      if(when_BankedScratchMemory_l242_65) begin
        banks_1_io_write_addr = _zz_io_write_addr_8;
      end
    end
    if(io_writeEn_9) begin
      if(when_BankedScratchMemory_l242_73) begin
        banks_1_io_write_addr = _zz_io_write_addr_9;
      end
    end
    if(io_writeEn_10) begin
      if(when_BankedScratchMemory_l242_81) begin
        banks_1_io_write_addr = _zz_io_write_addr_10;
      end
    end
    if(io_writeEn_11) begin
      if(when_BankedScratchMemory_l242_89) begin
        banks_1_io_write_addr = _zz_io_write_addr_11;
      end
    end
    if(io_writeEn_12) begin
      if(when_BankedScratchMemory_l242_97) begin
        banks_1_io_write_addr = _zz_io_write_addr_12;
      end
    end
    if(io_writeEn_13) begin
      if(when_BankedScratchMemory_l242_105) begin
        banks_1_io_write_addr = _zz_io_write_addr_13;
      end
    end
    if(io_writeEn_14) begin
      if(when_BankedScratchMemory_l242_113) begin
        banks_1_io_write_addr = _zz_io_write_addr_14;
      end
    end
    if(io_writeEn_15) begin
      if(when_BankedScratchMemory_l242_121) begin
        banks_1_io_write_addr = _zz_io_write_addr_15;
      end
    end
    if(io_writeEn_16) begin
      if(when_BankedScratchMemory_l242_129) begin
        banks_1_io_write_addr = _zz_io_write_addr_16;
      end
    end
    if(io_writeEn_17) begin
      if(when_BankedScratchMemory_l242_137) begin
        banks_1_io_write_addr = _zz_io_write_addr_17;
      end
    end
    if(io_writeEn_18) begin
      if(when_BankedScratchMemory_l242_145) begin
        banks_1_io_write_addr = _zz_io_write_addr_18;
      end
    end
    if(io_writeEn_19) begin
      if(when_BankedScratchMemory_l242_153) begin
        banks_1_io_write_addr = _zz_io_write_addr_19;
      end
    end
    if(io_writeEn_20) begin
      if(when_BankedScratchMemory_l242_161) begin
        banks_1_io_write_addr = _zz_io_write_addr_20;
      end
    end
    if(io_writeEn_21) begin
      if(when_BankedScratchMemory_l242_169) begin
        banks_1_io_write_addr = _zz_io_write_addr_21;
      end
    end
    if(io_writeEn_22) begin
      if(when_BankedScratchMemory_l242_177) begin
        banks_1_io_write_addr = _zz_io_write_addr_22;
      end
    end
    if(io_writeEn_23) begin
      if(when_BankedScratchMemory_l242_185) begin
        banks_1_io_write_addr = _zz_io_write_addr_23;
      end
    end
    if(io_writeEn_24) begin
      if(when_BankedScratchMemory_l242_193) begin
        banks_1_io_write_addr = _zz_io_write_addr_24;
      end
    end
    if(io_writeEn_25) begin
      if(when_BankedScratchMemory_l242_201) begin
        banks_1_io_write_addr = _zz_io_write_addr_25;
      end
    end
    if(io_writeEn_26) begin
      if(when_BankedScratchMemory_l242_209) begin
        banks_1_io_write_addr = _zz_io_write_addr_26;
      end
    end
    if(io_writeEn_27) begin
      if(when_BankedScratchMemory_l242_217) begin
        banks_1_io_write_addr = _zz_io_write_addr_27;
      end
    end
  end

  always @(*) begin
    banks_1_io_write_data = 32'h0;
    if(io_writeEn_0) begin
      if(when_BankedScratchMemory_l242_1) begin
        banks_1_io_write_data = io_writeData_0;
      end
    end
    if(io_writeEn_1) begin
      if(when_BankedScratchMemory_l242_9) begin
        banks_1_io_write_data = io_writeData_1;
      end
    end
    if(io_writeEn_2) begin
      if(when_BankedScratchMemory_l242_17) begin
        banks_1_io_write_data = io_writeData_2;
      end
    end
    if(io_writeEn_3) begin
      if(when_BankedScratchMemory_l242_25) begin
        banks_1_io_write_data = io_writeData_3;
      end
    end
    if(io_writeEn_4) begin
      if(when_BankedScratchMemory_l242_33) begin
        banks_1_io_write_data = io_writeData_4;
      end
    end
    if(io_writeEn_5) begin
      if(when_BankedScratchMemory_l242_41) begin
        banks_1_io_write_data = io_writeData_5;
      end
    end
    if(io_writeEn_6) begin
      if(when_BankedScratchMemory_l242_49) begin
        banks_1_io_write_data = io_writeData_6;
      end
    end
    if(io_writeEn_7) begin
      if(when_BankedScratchMemory_l242_57) begin
        banks_1_io_write_data = io_writeData_7;
      end
    end
    if(io_writeEn_8) begin
      if(when_BankedScratchMemory_l242_65) begin
        banks_1_io_write_data = io_writeData_8;
      end
    end
    if(io_writeEn_9) begin
      if(when_BankedScratchMemory_l242_73) begin
        banks_1_io_write_data = io_writeData_9;
      end
    end
    if(io_writeEn_10) begin
      if(when_BankedScratchMemory_l242_81) begin
        banks_1_io_write_data = io_writeData_10;
      end
    end
    if(io_writeEn_11) begin
      if(when_BankedScratchMemory_l242_89) begin
        banks_1_io_write_data = io_writeData_11;
      end
    end
    if(io_writeEn_12) begin
      if(when_BankedScratchMemory_l242_97) begin
        banks_1_io_write_data = io_writeData_12;
      end
    end
    if(io_writeEn_13) begin
      if(when_BankedScratchMemory_l242_105) begin
        banks_1_io_write_data = io_writeData_13;
      end
    end
    if(io_writeEn_14) begin
      if(when_BankedScratchMemory_l242_113) begin
        banks_1_io_write_data = io_writeData_14;
      end
    end
    if(io_writeEn_15) begin
      if(when_BankedScratchMemory_l242_121) begin
        banks_1_io_write_data = io_writeData_15;
      end
    end
    if(io_writeEn_16) begin
      if(when_BankedScratchMemory_l242_129) begin
        banks_1_io_write_data = io_writeData_16;
      end
    end
    if(io_writeEn_17) begin
      if(when_BankedScratchMemory_l242_137) begin
        banks_1_io_write_data = io_writeData_17;
      end
    end
    if(io_writeEn_18) begin
      if(when_BankedScratchMemory_l242_145) begin
        banks_1_io_write_data = io_writeData_18;
      end
    end
    if(io_writeEn_19) begin
      if(when_BankedScratchMemory_l242_153) begin
        banks_1_io_write_data = io_writeData_19;
      end
    end
    if(io_writeEn_20) begin
      if(when_BankedScratchMemory_l242_161) begin
        banks_1_io_write_data = io_writeData_20;
      end
    end
    if(io_writeEn_21) begin
      if(when_BankedScratchMemory_l242_169) begin
        banks_1_io_write_data = io_writeData_21;
      end
    end
    if(io_writeEn_22) begin
      if(when_BankedScratchMemory_l242_177) begin
        banks_1_io_write_data = io_writeData_22;
      end
    end
    if(io_writeEn_23) begin
      if(when_BankedScratchMemory_l242_185) begin
        banks_1_io_write_data = io_writeData_23;
      end
    end
    if(io_writeEn_24) begin
      if(when_BankedScratchMemory_l242_193) begin
        banks_1_io_write_data = io_writeData_24;
      end
    end
    if(io_writeEn_25) begin
      if(when_BankedScratchMemory_l242_201) begin
        banks_1_io_write_data = io_writeData_25;
      end
    end
    if(io_writeEn_26) begin
      if(when_BankedScratchMemory_l242_209) begin
        banks_1_io_write_data = io_writeData_26;
      end
    end
    if(io_writeEn_27) begin
      if(when_BankedScratchMemory_l242_217) begin
        banks_1_io_write_data = io_writeData_27;
      end
    end
  end

  always @(*) begin
    banks_2_io_write_en = 1'b0;
    if(io_writeEn_0) begin
      if(when_BankedScratchMemory_l242_2) begin
        banks_2_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_1) begin
      if(when_BankedScratchMemory_l242_10) begin
        banks_2_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_2) begin
      if(when_BankedScratchMemory_l242_18) begin
        banks_2_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_3) begin
      if(when_BankedScratchMemory_l242_26) begin
        banks_2_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_4) begin
      if(when_BankedScratchMemory_l242_34) begin
        banks_2_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_5) begin
      if(when_BankedScratchMemory_l242_42) begin
        banks_2_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_6) begin
      if(when_BankedScratchMemory_l242_50) begin
        banks_2_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_7) begin
      if(when_BankedScratchMemory_l242_58) begin
        banks_2_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_8) begin
      if(when_BankedScratchMemory_l242_66) begin
        banks_2_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_9) begin
      if(when_BankedScratchMemory_l242_74) begin
        banks_2_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_10) begin
      if(when_BankedScratchMemory_l242_82) begin
        banks_2_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_11) begin
      if(when_BankedScratchMemory_l242_90) begin
        banks_2_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_12) begin
      if(when_BankedScratchMemory_l242_98) begin
        banks_2_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_13) begin
      if(when_BankedScratchMemory_l242_106) begin
        banks_2_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_14) begin
      if(when_BankedScratchMemory_l242_114) begin
        banks_2_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_15) begin
      if(when_BankedScratchMemory_l242_122) begin
        banks_2_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_16) begin
      if(when_BankedScratchMemory_l242_130) begin
        banks_2_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_17) begin
      if(when_BankedScratchMemory_l242_138) begin
        banks_2_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_18) begin
      if(when_BankedScratchMemory_l242_146) begin
        banks_2_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_19) begin
      if(when_BankedScratchMemory_l242_154) begin
        banks_2_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_20) begin
      if(when_BankedScratchMemory_l242_162) begin
        banks_2_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_21) begin
      if(when_BankedScratchMemory_l242_170) begin
        banks_2_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_22) begin
      if(when_BankedScratchMemory_l242_178) begin
        banks_2_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_23) begin
      if(when_BankedScratchMemory_l242_186) begin
        banks_2_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_24) begin
      if(when_BankedScratchMemory_l242_194) begin
        banks_2_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_25) begin
      if(when_BankedScratchMemory_l242_202) begin
        banks_2_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_26) begin
      if(when_BankedScratchMemory_l242_210) begin
        banks_2_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_27) begin
      if(when_BankedScratchMemory_l242_218) begin
        banks_2_io_write_en = 1'b1;
      end
    end
  end

  always @(*) begin
    banks_2_io_write_addr = 8'h0;
    if(io_writeEn_0) begin
      if(when_BankedScratchMemory_l242_2) begin
        banks_2_io_write_addr = _zz_io_write_addr;
      end
    end
    if(io_writeEn_1) begin
      if(when_BankedScratchMemory_l242_10) begin
        banks_2_io_write_addr = _zz_io_write_addr_1;
      end
    end
    if(io_writeEn_2) begin
      if(when_BankedScratchMemory_l242_18) begin
        banks_2_io_write_addr = _zz_io_write_addr_2;
      end
    end
    if(io_writeEn_3) begin
      if(when_BankedScratchMemory_l242_26) begin
        banks_2_io_write_addr = _zz_io_write_addr_3;
      end
    end
    if(io_writeEn_4) begin
      if(when_BankedScratchMemory_l242_34) begin
        banks_2_io_write_addr = _zz_io_write_addr_4;
      end
    end
    if(io_writeEn_5) begin
      if(when_BankedScratchMemory_l242_42) begin
        banks_2_io_write_addr = _zz_io_write_addr_5;
      end
    end
    if(io_writeEn_6) begin
      if(when_BankedScratchMemory_l242_50) begin
        banks_2_io_write_addr = _zz_io_write_addr_6;
      end
    end
    if(io_writeEn_7) begin
      if(when_BankedScratchMemory_l242_58) begin
        banks_2_io_write_addr = _zz_io_write_addr_7;
      end
    end
    if(io_writeEn_8) begin
      if(when_BankedScratchMemory_l242_66) begin
        banks_2_io_write_addr = _zz_io_write_addr_8;
      end
    end
    if(io_writeEn_9) begin
      if(when_BankedScratchMemory_l242_74) begin
        banks_2_io_write_addr = _zz_io_write_addr_9;
      end
    end
    if(io_writeEn_10) begin
      if(when_BankedScratchMemory_l242_82) begin
        banks_2_io_write_addr = _zz_io_write_addr_10;
      end
    end
    if(io_writeEn_11) begin
      if(when_BankedScratchMemory_l242_90) begin
        banks_2_io_write_addr = _zz_io_write_addr_11;
      end
    end
    if(io_writeEn_12) begin
      if(when_BankedScratchMemory_l242_98) begin
        banks_2_io_write_addr = _zz_io_write_addr_12;
      end
    end
    if(io_writeEn_13) begin
      if(when_BankedScratchMemory_l242_106) begin
        banks_2_io_write_addr = _zz_io_write_addr_13;
      end
    end
    if(io_writeEn_14) begin
      if(when_BankedScratchMemory_l242_114) begin
        banks_2_io_write_addr = _zz_io_write_addr_14;
      end
    end
    if(io_writeEn_15) begin
      if(when_BankedScratchMemory_l242_122) begin
        banks_2_io_write_addr = _zz_io_write_addr_15;
      end
    end
    if(io_writeEn_16) begin
      if(when_BankedScratchMemory_l242_130) begin
        banks_2_io_write_addr = _zz_io_write_addr_16;
      end
    end
    if(io_writeEn_17) begin
      if(when_BankedScratchMemory_l242_138) begin
        banks_2_io_write_addr = _zz_io_write_addr_17;
      end
    end
    if(io_writeEn_18) begin
      if(when_BankedScratchMemory_l242_146) begin
        banks_2_io_write_addr = _zz_io_write_addr_18;
      end
    end
    if(io_writeEn_19) begin
      if(when_BankedScratchMemory_l242_154) begin
        banks_2_io_write_addr = _zz_io_write_addr_19;
      end
    end
    if(io_writeEn_20) begin
      if(when_BankedScratchMemory_l242_162) begin
        banks_2_io_write_addr = _zz_io_write_addr_20;
      end
    end
    if(io_writeEn_21) begin
      if(when_BankedScratchMemory_l242_170) begin
        banks_2_io_write_addr = _zz_io_write_addr_21;
      end
    end
    if(io_writeEn_22) begin
      if(when_BankedScratchMemory_l242_178) begin
        banks_2_io_write_addr = _zz_io_write_addr_22;
      end
    end
    if(io_writeEn_23) begin
      if(when_BankedScratchMemory_l242_186) begin
        banks_2_io_write_addr = _zz_io_write_addr_23;
      end
    end
    if(io_writeEn_24) begin
      if(when_BankedScratchMemory_l242_194) begin
        banks_2_io_write_addr = _zz_io_write_addr_24;
      end
    end
    if(io_writeEn_25) begin
      if(when_BankedScratchMemory_l242_202) begin
        banks_2_io_write_addr = _zz_io_write_addr_25;
      end
    end
    if(io_writeEn_26) begin
      if(when_BankedScratchMemory_l242_210) begin
        banks_2_io_write_addr = _zz_io_write_addr_26;
      end
    end
    if(io_writeEn_27) begin
      if(when_BankedScratchMemory_l242_218) begin
        banks_2_io_write_addr = _zz_io_write_addr_27;
      end
    end
  end

  always @(*) begin
    banks_2_io_write_data = 32'h0;
    if(io_writeEn_0) begin
      if(when_BankedScratchMemory_l242_2) begin
        banks_2_io_write_data = io_writeData_0;
      end
    end
    if(io_writeEn_1) begin
      if(when_BankedScratchMemory_l242_10) begin
        banks_2_io_write_data = io_writeData_1;
      end
    end
    if(io_writeEn_2) begin
      if(when_BankedScratchMemory_l242_18) begin
        banks_2_io_write_data = io_writeData_2;
      end
    end
    if(io_writeEn_3) begin
      if(when_BankedScratchMemory_l242_26) begin
        banks_2_io_write_data = io_writeData_3;
      end
    end
    if(io_writeEn_4) begin
      if(when_BankedScratchMemory_l242_34) begin
        banks_2_io_write_data = io_writeData_4;
      end
    end
    if(io_writeEn_5) begin
      if(when_BankedScratchMemory_l242_42) begin
        banks_2_io_write_data = io_writeData_5;
      end
    end
    if(io_writeEn_6) begin
      if(when_BankedScratchMemory_l242_50) begin
        banks_2_io_write_data = io_writeData_6;
      end
    end
    if(io_writeEn_7) begin
      if(when_BankedScratchMemory_l242_58) begin
        banks_2_io_write_data = io_writeData_7;
      end
    end
    if(io_writeEn_8) begin
      if(when_BankedScratchMemory_l242_66) begin
        banks_2_io_write_data = io_writeData_8;
      end
    end
    if(io_writeEn_9) begin
      if(when_BankedScratchMemory_l242_74) begin
        banks_2_io_write_data = io_writeData_9;
      end
    end
    if(io_writeEn_10) begin
      if(when_BankedScratchMemory_l242_82) begin
        banks_2_io_write_data = io_writeData_10;
      end
    end
    if(io_writeEn_11) begin
      if(when_BankedScratchMemory_l242_90) begin
        banks_2_io_write_data = io_writeData_11;
      end
    end
    if(io_writeEn_12) begin
      if(when_BankedScratchMemory_l242_98) begin
        banks_2_io_write_data = io_writeData_12;
      end
    end
    if(io_writeEn_13) begin
      if(when_BankedScratchMemory_l242_106) begin
        banks_2_io_write_data = io_writeData_13;
      end
    end
    if(io_writeEn_14) begin
      if(when_BankedScratchMemory_l242_114) begin
        banks_2_io_write_data = io_writeData_14;
      end
    end
    if(io_writeEn_15) begin
      if(when_BankedScratchMemory_l242_122) begin
        banks_2_io_write_data = io_writeData_15;
      end
    end
    if(io_writeEn_16) begin
      if(when_BankedScratchMemory_l242_130) begin
        banks_2_io_write_data = io_writeData_16;
      end
    end
    if(io_writeEn_17) begin
      if(when_BankedScratchMemory_l242_138) begin
        banks_2_io_write_data = io_writeData_17;
      end
    end
    if(io_writeEn_18) begin
      if(when_BankedScratchMemory_l242_146) begin
        banks_2_io_write_data = io_writeData_18;
      end
    end
    if(io_writeEn_19) begin
      if(when_BankedScratchMemory_l242_154) begin
        banks_2_io_write_data = io_writeData_19;
      end
    end
    if(io_writeEn_20) begin
      if(when_BankedScratchMemory_l242_162) begin
        banks_2_io_write_data = io_writeData_20;
      end
    end
    if(io_writeEn_21) begin
      if(when_BankedScratchMemory_l242_170) begin
        banks_2_io_write_data = io_writeData_21;
      end
    end
    if(io_writeEn_22) begin
      if(when_BankedScratchMemory_l242_178) begin
        banks_2_io_write_data = io_writeData_22;
      end
    end
    if(io_writeEn_23) begin
      if(when_BankedScratchMemory_l242_186) begin
        banks_2_io_write_data = io_writeData_23;
      end
    end
    if(io_writeEn_24) begin
      if(when_BankedScratchMemory_l242_194) begin
        banks_2_io_write_data = io_writeData_24;
      end
    end
    if(io_writeEn_25) begin
      if(when_BankedScratchMemory_l242_202) begin
        banks_2_io_write_data = io_writeData_25;
      end
    end
    if(io_writeEn_26) begin
      if(when_BankedScratchMemory_l242_210) begin
        banks_2_io_write_data = io_writeData_26;
      end
    end
    if(io_writeEn_27) begin
      if(when_BankedScratchMemory_l242_218) begin
        banks_2_io_write_data = io_writeData_27;
      end
    end
  end

  always @(*) begin
    banks_3_io_write_en = 1'b0;
    if(io_writeEn_0) begin
      if(when_BankedScratchMemory_l242_3) begin
        banks_3_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_1) begin
      if(when_BankedScratchMemory_l242_11) begin
        banks_3_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_2) begin
      if(when_BankedScratchMemory_l242_19) begin
        banks_3_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_3) begin
      if(when_BankedScratchMemory_l242_27) begin
        banks_3_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_4) begin
      if(when_BankedScratchMemory_l242_35) begin
        banks_3_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_5) begin
      if(when_BankedScratchMemory_l242_43) begin
        banks_3_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_6) begin
      if(when_BankedScratchMemory_l242_51) begin
        banks_3_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_7) begin
      if(when_BankedScratchMemory_l242_59) begin
        banks_3_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_8) begin
      if(when_BankedScratchMemory_l242_67) begin
        banks_3_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_9) begin
      if(when_BankedScratchMemory_l242_75) begin
        banks_3_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_10) begin
      if(when_BankedScratchMemory_l242_83) begin
        banks_3_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_11) begin
      if(when_BankedScratchMemory_l242_91) begin
        banks_3_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_12) begin
      if(when_BankedScratchMemory_l242_99) begin
        banks_3_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_13) begin
      if(when_BankedScratchMemory_l242_107) begin
        banks_3_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_14) begin
      if(when_BankedScratchMemory_l242_115) begin
        banks_3_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_15) begin
      if(when_BankedScratchMemory_l242_123) begin
        banks_3_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_16) begin
      if(when_BankedScratchMemory_l242_131) begin
        banks_3_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_17) begin
      if(when_BankedScratchMemory_l242_139) begin
        banks_3_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_18) begin
      if(when_BankedScratchMemory_l242_147) begin
        banks_3_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_19) begin
      if(when_BankedScratchMemory_l242_155) begin
        banks_3_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_20) begin
      if(when_BankedScratchMemory_l242_163) begin
        banks_3_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_21) begin
      if(when_BankedScratchMemory_l242_171) begin
        banks_3_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_22) begin
      if(when_BankedScratchMemory_l242_179) begin
        banks_3_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_23) begin
      if(when_BankedScratchMemory_l242_187) begin
        banks_3_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_24) begin
      if(when_BankedScratchMemory_l242_195) begin
        banks_3_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_25) begin
      if(when_BankedScratchMemory_l242_203) begin
        banks_3_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_26) begin
      if(when_BankedScratchMemory_l242_211) begin
        banks_3_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_27) begin
      if(when_BankedScratchMemory_l242_219) begin
        banks_3_io_write_en = 1'b1;
      end
    end
  end

  always @(*) begin
    banks_3_io_write_addr = 8'h0;
    if(io_writeEn_0) begin
      if(when_BankedScratchMemory_l242_3) begin
        banks_3_io_write_addr = _zz_io_write_addr;
      end
    end
    if(io_writeEn_1) begin
      if(when_BankedScratchMemory_l242_11) begin
        banks_3_io_write_addr = _zz_io_write_addr_1;
      end
    end
    if(io_writeEn_2) begin
      if(when_BankedScratchMemory_l242_19) begin
        banks_3_io_write_addr = _zz_io_write_addr_2;
      end
    end
    if(io_writeEn_3) begin
      if(when_BankedScratchMemory_l242_27) begin
        banks_3_io_write_addr = _zz_io_write_addr_3;
      end
    end
    if(io_writeEn_4) begin
      if(when_BankedScratchMemory_l242_35) begin
        banks_3_io_write_addr = _zz_io_write_addr_4;
      end
    end
    if(io_writeEn_5) begin
      if(when_BankedScratchMemory_l242_43) begin
        banks_3_io_write_addr = _zz_io_write_addr_5;
      end
    end
    if(io_writeEn_6) begin
      if(when_BankedScratchMemory_l242_51) begin
        banks_3_io_write_addr = _zz_io_write_addr_6;
      end
    end
    if(io_writeEn_7) begin
      if(when_BankedScratchMemory_l242_59) begin
        banks_3_io_write_addr = _zz_io_write_addr_7;
      end
    end
    if(io_writeEn_8) begin
      if(when_BankedScratchMemory_l242_67) begin
        banks_3_io_write_addr = _zz_io_write_addr_8;
      end
    end
    if(io_writeEn_9) begin
      if(when_BankedScratchMemory_l242_75) begin
        banks_3_io_write_addr = _zz_io_write_addr_9;
      end
    end
    if(io_writeEn_10) begin
      if(when_BankedScratchMemory_l242_83) begin
        banks_3_io_write_addr = _zz_io_write_addr_10;
      end
    end
    if(io_writeEn_11) begin
      if(when_BankedScratchMemory_l242_91) begin
        banks_3_io_write_addr = _zz_io_write_addr_11;
      end
    end
    if(io_writeEn_12) begin
      if(when_BankedScratchMemory_l242_99) begin
        banks_3_io_write_addr = _zz_io_write_addr_12;
      end
    end
    if(io_writeEn_13) begin
      if(when_BankedScratchMemory_l242_107) begin
        banks_3_io_write_addr = _zz_io_write_addr_13;
      end
    end
    if(io_writeEn_14) begin
      if(when_BankedScratchMemory_l242_115) begin
        banks_3_io_write_addr = _zz_io_write_addr_14;
      end
    end
    if(io_writeEn_15) begin
      if(when_BankedScratchMemory_l242_123) begin
        banks_3_io_write_addr = _zz_io_write_addr_15;
      end
    end
    if(io_writeEn_16) begin
      if(when_BankedScratchMemory_l242_131) begin
        banks_3_io_write_addr = _zz_io_write_addr_16;
      end
    end
    if(io_writeEn_17) begin
      if(when_BankedScratchMemory_l242_139) begin
        banks_3_io_write_addr = _zz_io_write_addr_17;
      end
    end
    if(io_writeEn_18) begin
      if(when_BankedScratchMemory_l242_147) begin
        banks_3_io_write_addr = _zz_io_write_addr_18;
      end
    end
    if(io_writeEn_19) begin
      if(when_BankedScratchMemory_l242_155) begin
        banks_3_io_write_addr = _zz_io_write_addr_19;
      end
    end
    if(io_writeEn_20) begin
      if(when_BankedScratchMemory_l242_163) begin
        banks_3_io_write_addr = _zz_io_write_addr_20;
      end
    end
    if(io_writeEn_21) begin
      if(when_BankedScratchMemory_l242_171) begin
        banks_3_io_write_addr = _zz_io_write_addr_21;
      end
    end
    if(io_writeEn_22) begin
      if(when_BankedScratchMemory_l242_179) begin
        banks_3_io_write_addr = _zz_io_write_addr_22;
      end
    end
    if(io_writeEn_23) begin
      if(when_BankedScratchMemory_l242_187) begin
        banks_3_io_write_addr = _zz_io_write_addr_23;
      end
    end
    if(io_writeEn_24) begin
      if(when_BankedScratchMemory_l242_195) begin
        banks_3_io_write_addr = _zz_io_write_addr_24;
      end
    end
    if(io_writeEn_25) begin
      if(when_BankedScratchMemory_l242_203) begin
        banks_3_io_write_addr = _zz_io_write_addr_25;
      end
    end
    if(io_writeEn_26) begin
      if(when_BankedScratchMemory_l242_211) begin
        banks_3_io_write_addr = _zz_io_write_addr_26;
      end
    end
    if(io_writeEn_27) begin
      if(when_BankedScratchMemory_l242_219) begin
        banks_3_io_write_addr = _zz_io_write_addr_27;
      end
    end
  end

  always @(*) begin
    banks_3_io_write_data = 32'h0;
    if(io_writeEn_0) begin
      if(when_BankedScratchMemory_l242_3) begin
        banks_3_io_write_data = io_writeData_0;
      end
    end
    if(io_writeEn_1) begin
      if(when_BankedScratchMemory_l242_11) begin
        banks_3_io_write_data = io_writeData_1;
      end
    end
    if(io_writeEn_2) begin
      if(when_BankedScratchMemory_l242_19) begin
        banks_3_io_write_data = io_writeData_2;
      end
    end
    if(io_writeEn_3) begin
      if(when_BankedScratchMemory_l242_27) begin
        banks_3_io_write_data = io_writeData_3;
      end
    end
    if(io_writeEn_4) begin
      if(when_BankedScratchMemory_l242_35) begin
        banks_3_io_write_data = io_writeData_4;
      end
    end
    if(io_writeEn_5) begin
      if(when_BankedScratchMemory_l242_43) begin
        banks_3_io_write_data = io_writeData_5;
      end
    end
    if(io_writeEn_6) begin
      if(when_BankedScratchMemory_l242_51) begin
        banks_3_io_write_data = io_writeData_6;
      end
    end
    if(io_writeEn_7) begin
      if(when_BankedScratchMemory_l242_59) begin
        banks_3_io_write_data = io_writeData_7;
      end
    end
    if(io_writeEn_8) begin
      if(when_BankedScratchMemory_l242_67) begin
        banks_3_io_write_data = io_writeData_8;
      end
    end
    if(io_writeEn_9) begin
      if(when_BankedScratchMemory_l242_75) begin
        banks_3_io_write_data = io_writeData_9;
      end
    end
    if(io_writeEn_10) begin
      if(when_BankedScratchMemory_l242_83) begin
        banks_3_io_write_data = io_writeData_10;
      end
    end
    if(io_writeEn_11) begin
      if(when_BankedScratchMemory_l242_91) begin
        banks_3_io_write_data = io_writeData_11;
      end
    end
    if(io_writeEn_12) begin
      if(when_BankedScratchMemory_l242_99) begin
        banks_3_io_write_data = io_writeData_12;
      end
    end
    if(io_writeEn_13) begin
      if(when_BankedScratchMemory_l242_107) begin
        banks_3_io_write_data = io_writeData_13;
      end
    end
    if(io_writeEn_14) begin
      if(when_BankedScratchMemory_l242_115) begin
        banks_3_io_write_data = io_writeData_14;
      end
    end
    if(io_writeEn_15) begin
      if(when_BankedScratchMemory_l242_123) begin
        banks_3_io_write_data = io_writeData_15;
      end
    end
    if(io_writeEn_16) begin
      if(when_BankedScratchMemory_l242_131) begin
        banks_3_io_write_data = io_writeData_16;
      end
    end
    if(io_writeEn_17) begin
      if(when_BankedScratchMemory_l242_139) begin
        banks_3_io_write_data = io_writeData_17;
      end
    end
    if(io_writeEn_18) begin
      if(when_BankedScratchMemory_l242_147) begin
        banks_3_io_write_data = io_writeData_18;
      end
    end
    if(io_writeEn_19) begin
      if(when_BankedScratchMemory_l242_155) begin
        banks_3_io_write_data = io_writeData_19;
      end
    end
    if(io_writeEn_20) begin
      if(when_BankedScratchMemory_l242_163) begin
        banks_3_io_write_data = io_writeData_20;
      end
    end
    if(io_writeEn_21) begin
      if(when_BankedScratchMemory_l242_171) begin
        banks_3_io_write_data = io_writeData_21;
      end
    end
    if(io_writeEn_22) begin
      if(when_BankedScratchMemory_l242_179) begin
        banks_3_io_write_data = io_writeData_22;
      end
    end
    if(io_writeEn_23) begin
      if(when_BankedScratchMemory_l242_187) begin
        banks_3_io_write_data = io_writeData_23;
      end
    end
    if(io_writeEn_24) begin
      if(when_BankedScratchMemory_l242_195) begin
        banks_3_io_write_data = io_writeData_24;
      end
    end
    if(io_writeEn_25) begin
      if(when_BankedScratchMemory_l242_203) begin
        banks_3_io_write_data = io_writeData_25;
      end
    end
    if(io_writeEn_26) begin
      if(when_BankedScratchMemory_l242_211) begin
        banks_3_io_write_data = io_writeData_26;
      end
    end
    if(io_writeEn_27) begin
      if(when_BankedScratchMemory_l242_219) begin
        banks_3_io_write_data = io_writeData_27;
      end
    end
  end

  always @(*) begin
    banks_4_io_write_en = 1'b0;
    if(io_writeEn_0) begin
      if(when_BankedScratchMemory_l242_4) begin
        banks_4_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_1) begin
      if(when_BankedScratchMemory_l242_12) begin
        banks_4_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_2) begin
      if(when_BankedScratchMemory_l242_20) begin
        banks_4_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_3) begin
      if(when_BankedScratchMemory_l242_28) begin
        banks_4_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_4) begin
      if(when_BankedScratchMemory_l242_36) begin
        banks_4_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_5) begin
      if(when_BankedScratchMemory_l242_44) begin
        banks_4_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_6) begin
      if(when_BankedScratchMemory_l242_52) begin
        banks_4_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_7) begin
      if(when_BankedScratchMemory_l242_60) begin
        banks_4_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_8) begin
      if(when_BankedScratchMemory_l242_68) begin
        banks_4_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_9) begin
      if(when_BankedScratchMemory_l242_76) begin
        banks_4_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_10) begin
      if(when_BankedScratchMemory_l242_84) begin
        banks_4_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_11) begin
      if(when_BankedScratchMemory_l242_92) begin
        banks_4_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_12) begin
      if(when_BankedScratchMemory_l242_100) begin
        banks_4_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_13) begin
      if(when_BankedScratchMemory_l242_108) begin
        banks_4_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_14) begin
      if(when_BankedScratchMemory_l242_116) begin
        banks_4_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_15) begin
      if(when_BankedScratchMemory_l242_124) begin
        banks_4_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_16) begin
      if(when_BankedScratchMemory_l242_132) begin
        banks_4_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_17) begin
      if(when_BankedScratchMemory_l242_140) begin
        banks_4_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_18) begin
      if(when_BankedScratchMemory_l242_148) begin
        banks_4_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_19) begin
      if(when_BankedScratchMemory_l242_156) begin
        banks_4_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_20) begin
      if(when_BankedScratchMemory_l242_164) begin
        banks_4_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_21) begin
      if(when_BankedScratchMemory_l242_172) begin
        banks_4_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_22) begin
      if(when_BankedScratchMemory_l242_180) begin
        banks_4_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_23) begin
      if(when_BankedScratchMemory_l242_188) begin
        banks_4_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_24) begin
      if(when_BankedScratchMemory_l242_196) begin
        banks_4_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_25) begin
      if(when_BankedScratchMemory_l242_204) begin
        banks_4_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_26) begin
      if(when_BankedScratchMemory_l242_212) begin
        banks_4_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_27) begin
      if(when_BankedScratchMemory_l242_220) begin
        banks_4_io_write_en = 1'b1;
      end
    end
  end

  always @(*) begin
    banks_4_io_write_addr = 8'h0;
    if(io_writeEn_0) begin
      if(when_BankedScratchMemory_l242_4) begin
        banks_4_io_write_addr = _zz_io_write_addr;
      end
    end
    if(io_writeEn_1) begin
      if(when_BankedScratchMemory_l242_12) begin
        banks_4_io_write_addr = _zz_io_write_addr_1;
      end
    end
    if(io_writeEn_2) begin
      if(when_BankedScratchMemory_l242_20) begin
        banks_4_io_write_addr = _zz_io_write_addr_2;
      end
    end
    if(io_writeEn_3) begin
      if(when_BankedScratchMemory_l242_28) begin
        banks_4_io_write_addr = _zz_io_write_addr_3;
      end
    end
    if(io_writeEn_4) begin
      if(when_BankedScratchMemory_l242_36) begin
        banks_4_io_write_addr = _zz_io_write_addr_4;
      end
    end
    if(io_writeEn_5) begin
      if(when_BankedScratchMemory_l242_44) begin
        banks_4_io_write_addr = _zz_io_write_addr_5;
      end
    end
    if(io_writeEn_6) begin
      if(when_BankedScratchMemory_l242_52) begin
        banks_4_io_write_addr = _zz_io_write_addr_6;
      end
    end
    if(io_writeEn_7) begin
      if(when_BankedScratchMemory_l242_60) begin
        banks_4_io_write_addr = _zz_io_write_addr_7;
      end
    end
    if(io_writeEn_8) begin
      if(when_BankedScratchMemory_l242_68) begin
        banks_4_io_write_addr = _zz_io_write_addr_8;
      end
    end
    if(io_writeEn_9) begin
      if(when_BankedScratchMemory_l242_76) begin
        banks_4_io_write_addr = _zz_io_write_addr_9;
      end
    end
    if(io_writeEn_10) begin
      if(when_BankedScratchMemory_l242_84) begin
        banks_4_io_write_addr = _zz_io_write_addr_10;
      end
    end
    if(io_writeEn_11) begin
      if(when_BankedScratchMemory_l242_92) begin
        banks_4_io_write_addr = _zz_io_write_addr_11;
      end
    end
    if(io_writeEn_12) begin
      if(when_BankedScratchMemory_l242_100) begin
        banks_4_io_write_addr = _zz_io_write_addr_12;
      end
    end
    if(io_writeEn_13) begin
      if(when_BankedScratchMemory_l242_108) begin
        banks_4_io_write_addr = _zz_io_write_addr_13;
      end
    end
    if(io_writeEn_14) begin
      if(when_BankedScratchMemory_l242_116) begin
        banks_4_io_write_addr = _zz_io_write_addr_14;
      end
    end
    if(io_writeEn_15) begin
      if(when_BankedScratchMemory_l242_124) begin
        banks_4_io_write_addr = _zz_io_write_addr_15;
      end
    end
    if(io_writeEn_16) begin
      if(when_BankedScratchMemory_l242_132) begin
        banks_4_io_write_addr = _zz_io_write_addr_16;
      end
    end
    if(io_writeEn_17) begin
      if(when_BankedScratchMemory_l242_140) begin
        banks_4_io_write_addr = _zz_io_write_addr_17;
      end
    end
    if(io_writeEn_18) begin
      if(when_BankedScratchMemory_l242_148) begin
        banks_4_io_write_addr = _zz_io_write_addr_18;
      end
    end
    if(io_writeEn_19) begin
      if(when_BankedScratchMemory_l242_156) begin
        banks_4_io_write_addr = _zz_io_write_addr_19;
      end
    end
    if(io_writeEn_20) begin
      if(when_BankedScratchMemory_l242_164) begin
        banks_4_io_write_addr = _zz_io_write_addr_20;
      end
    end
    if(io_writeEn_21) begin
      if(when_BankedScratchMemory_l242_172) begin
        banks_4_io_write_addr = _zz_io_write_addr_21;
      end
    end
    if(io_writeEn_22) begin
      if(when_BankedScratchMemory_l242_180) begin
        banks_4_io_write_addr = _zz_io_write_addr_22;
      end
    end
    if(io_writeEn_23) begin
      if(when_BankedScratchMemory_l242_188) begin
        banks_4_io_write_addr = _zz_io_write_addr_23;
      end
    end
    if(io_writeEn_24) begin
      if(when_BankedScratchMemory_l242_196) begin
        banks_4_io_write_addr = _zz_io_write_addr_24;
      end
    end
    if(io_writeEn_25) begin
      if(when_BankedScratchMemory_l242_204) begin
        banks_4_io_write_addr = _zz_io_write_addr_25;
      end
    end
    if(io_writeEn_26) begin
      if(when_BankedScratchMemory_l242_212) begin
        banks_4_io_write_addr = _zz_io_write_addr_26;
      end
    end
    if(io_writeEn_27) begin
      if(when_BankedScratchMemory_l242_220) begin
        banks_4_io_write_addr = _zz_io_write_addr_27;
      end
    end
  end

  always @(*) begin
    banks_4_io_write_data = 32'h0;
    if(io_writeEn_0) begin
      if(when_BankedScratchMemory_l242_4) begin
        banks_4_io_write_data = io_writeData_0;
      end
    end
    if(io_writeEn_1) begin
      if(when_BankedScratchMemory_l242_12) begin
        banks_4_io_write_data = io_writeData_1;
      end
    end
    if(io_writeEn_2) begin
      if(when_BankedScratchMemory_l242_20) begin
        banks_4_io_write_data = io_writeData_2;
      end
    end
    if(io_writeEn_3) begin
      if(when_BankedScratchMemory_l242_28) begin
        banks_4_io_write_data = io_writeData_3;
      end
    end
    if(io_writeEn_4) begin
      if(when_BankedScratchMemory_l242_36) begin
        banks_4_io_write_data = io_writeData_4;
      end
    end
    if(io_writeEn_5) begin
      if(when_BankedScratchMemory_l242_44) begin
        banks_4_io_write_data = io_writeData_5;
      end
    end
    if(io_writeEn_6) begin
      if(when_BankedScratchMemory_l242_52) begin
        banks_4_io_write_data = io_writeData_6;
      end
    end
    if(io_writeEn_7) begin
      if(when_BankedScratchMemory_l242_60) begin
        banks_4_io_write_data = io_writeData_7;
      end
    end
    if(io_writeEn_8) begin
      if(when_BankedScratchMemory_l242_68) begin
        banks_4_io_write_data = io_writeData_8;
      end
    end
    if(io_writeEn_9) begin
      if(when_BankedScratchMemory_l242_76) begin
        banks_4_io_write_data = io_writeData_9;
      end
    end
    if(io_writeEn_10) begin
      if(when_BankedScratchMemory_l242_84) begin
        banks_4_io_write_data = io_writeData_10;
      end
    end
    if(io_writeEn_11) begin
      if(when_BankedScratchMemory_l242_92) begin
        banks_4_io_write_data = io_writeData_11;
      end
    end
    if(io_writeEn_12) begin
      if(when_BankedScratchMemory_l242_100) begin
        banks_4_io_write_data = io_writeData_12;
      end
    end
    if(io_writeEn_13) begin
      if(when_BankedScratchMemory_l242_108) begin
        banks_4_io_write_data = io_writeData_13;
      end
    end
    if(io_writeEn_14) begin
      if(when_BankedScratchMemory_l242_116) begin
        banks_4_io_write_data = io_writeData_14;
      end
    end
    if(io_writeEn_15) begin
      if(when_BankedScratchMemory_l242_124) begin
        banks_4_io_write_data = io_writeData_15;
      end
    end
    if(io_writeEn_16) begin
      if(when_BankedScratchMemory_l242_132) begin
        banks_4_io_write_data = io_writeData_16;
      end
    end
    if(io_writeEn_17) begin
      if(when_BankedScratchMemory_l242_140) begin
        banks_4_io_write_data = io_writeData_17;
      end
    end
    if(io_writeEn_18) begin
      if(when_BankedScratchMemory_l242_148) begin
        banks_4_io_write_data = io_writeData_18;
      end
    end
    if(io_writeEn_19) begin
      if(when_BankedScratchMemory_l242_156) begin
        banks_4_io_write_data = io_writeData_19;
      end
    end
    if(io_writeEn_20) begin
      if(when_BankedScratchMemory_l242_164) begin
        banks_4_io_write_data = io_writeData_20;
      end
    end
    if(io_writeEn_21) begin
      if(when_BankedScratchMemory_l242_172) begin
        banks_4_io_write_data = io_writeData_21;
      end
    end
    if(io_writeEn_22) begin
      if(when_BankedScratchMemory_l242_180) begin
        banks_4_io_write_data = io_writeData_22;
      end
    end
    if(io_writeEn_23) begin
      if(when_BankedScratchMemory_l242_188) begin
        banks_4_io_write_data = io_writeData_23;
      end
    end
    if(io_writeEn_24) begin
      if(when_BankedScratchMemory_l242_196) begin
        banks_4_io_write_data = io_writeData_24;
      end
    end
    if(io_writeEn_25) begin
      if(when_BankedScratchMemory_l242_204) begin
        banks_4_io_write_data = io_writeData_25;
      end
    end
    if(io_writeEn_26) begin
      if(when_BankedScratchMemory_l242_212) begin
        banks_4_io_write_data = io_writeData_26;
      end
    end
    if(io_writeEn_27) begin
      if(when_BankedScratchMemory_l242_220) begin
        banks_4_io_write_data = io_writeData_27;
      end
    end
  end

  always @(*) begin
    banks_5_io_write_en = 1'b0;
    if(io_writeEn_0) begin
      if(when_BankedScratchMemory_l242_5) begin
        banks_5_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_1) begin
      if(when_BankedScratchMemory_l242_13) begin
        banks_5_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_2) begin
      if(when_BankedScratchMemory_l242_21) begin
        banks_5_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_3) begin
      if(when_BankedScratchMemory_l242_29) begin
        banks_5_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_4) begin
      if(when_BankedScratchMemory_l242_37) begin
        banks_5_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_5) begin
      if(when_BankedScratchMemory_l242_45) begin
        banks_5_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_6) begin
      if(when_BankedScratchMemory_l242_53) begin
        banks_5_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_7) begin
      if(when_BankedScratchMemory_l242_61) begin
        banks_5_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_8) begin
      if(when_BankedScratchMemory_l242_69) begin
        banks_5_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_9) begin
      if(when_BankedScratchMemory_l242_77) begin
        banks_5_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_10) begin
      if(when_BankedScratchMemory_l242_85) begin
        banks_5_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_11) begin
      if(when_BankedScratchMemory_l242_93) begin
        banks_5_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_12) begin
      if(when_BankedScratchMemory_l242_101) begin
        banks_5_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_13) begin
      if(when_BankedScratchMemory_l242_109) begin
        banks_5_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_14) begin
      if(when_BankedScratchMemory_l242_117) begin
        banks_5_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_15) begin
      if(when_BankedScratchMemory_l242_125) begin
        banks_5_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_16) begin
      if(when_BankedScratchMemory_l242_133) begin
        banks_5_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_17) begin
      if(when_BankedScratchMemory_l242_141) begin
        banks_5_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_18) begin
      if(when_BankedScratchMemory_l242_149) begin
        banks_5_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_19) begin
      if(when_BankedScratchMemory_l242_157) begin
        banks_5_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_20) begin
      if(when_BankedScratchMemory_l242_165) begin
        banks_5_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_21) begin
      if(when_BankedScratchMemory_l242_173) begin
        banks_5_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_22) begin
      if(when_BankedScratchMemory_l242_181) begin
        banks_5_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_23) begin
      if(when_BankedScratchMemory_l242_189) begin
        banks_5_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_24) begin
      if(when_BankedScratchMemory_l242_197) begin
        banks_5_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_25) begin
      if(when_BankedScratchMemory_l242_205) begin
        banks_5_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_26) begin
      if(when_BankedScratchMemory_l242_213) begin
        banks_5_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_27) begin
      if(when_BankedScratchMemory_l242_221) begin
        banks_5_io_write_en = 1'b1;
      end
    end
  end

  always @(*) begin
    banks_5_io_write_addr = 8'h0;
    if(io_writeEn_0) begin
      if(when_BankedScratchMemory_l242_5) begin
        banks_5_io_write_addr = _zz_io_write_addr;
      end
    end
    if(io_writeEn_1) begin
      if(when_BankedScratchMemory_l242_13) begin
        banks_5_io_write_addr = _zz_io_write_addr_1;
      end
    end
    if(io_writeEn_2) begin
      if(when_BankedScratchMemory_l242_21) begin
        banks_5_io_write_addr = _zz_io_write_addr_2;
      end
    end
    if(io_writeEn_3) begin
      if(when_BankedScratchMemory_l242_29) begin
        banks_5_io_write_addr = _zz_io_write_addr_3;
      end
    end
    if(io_writeEn_4) begin
      if(when_BankedScratchMemory_l242_37) begin
        banks_5_io_write_addr = _zz_io_write_addr_4;
      end
    end
    if(io_writeEn_5) begin
      if(when_BankedScratchMemory_l242_45) begin
        banks_5_io_write_addr = _zz_io_write_addr_5;
      end
    end
    if(io_writeEn_6) begin
      if(when_BankedScratchMemory_l242_53) begin
        banks_5_io_write_addr = _zz_io_write_addr_6;
      end
    end
    if(io_writeEn_7) begin
      if(when_BankedScratchMemory_l242_61) begin
        banks_5_io_write_addr = _zz_io_write_addr_7;
      end
    end
    if(io_writeEn_8) begin
      if(when_BankedScratchMemory_l242_69) begin
        banks_5_io_write_addr = _zz_io_write_addr_8;
      end
    end
    if(io_writeEn_9) begin
      if(when_BankedScratchMemory_l242_77) begin
        banks_5_io_write_addr = _zz_io_write_addr_9;
      end
    end
    if(io_writeEn_10) begin
      if(when_BankedScratchMemory_l242_85) begin
        banks_5_io_write_addr = _zz_io_write_addr_10;
      end
    end
    if(io_writeEn_11) begin
      if(when_BankedScratchMemory_l242_93) begin
        banks_5_io_write_addr = _zz_io_write_addr_11;
      end
    end
    if(io_writeEn_12) begin
      if(when_BankedScratchMemory_l242_101) begin
        banks_5_io_write_addr = _zz_io_write_addr_12;
      end
    end
    if(io_writeEn_13) begin
      if(when_BankedScratchMemory_l242_109) begin
        banks_5_io_write_addr = _zz_io_write_addr_13;
      end
    end
    if(io_writeEn_14) begin
      if(when_BankedScratchMemory_l242_117) begin
        banks_5_io_write_addr = _zz_io_write_addr_14;
      end
    end
    if(io_writeEn_15) begin
      if(when_BankedScratchMemory_l242_125) begin
        banks_5_io_write_addr = _zz_io_write_addr_15;
      end
    end
    if(io_writeEn_16) begin
      if(when_BankedScratchMemory_l242_133) begin
        banks_5_io_write_addr = _zz_io_write_addr_16;
      end
    end
    if(io_writeEn_17) begin
      if(when_BankedScratchMemory_l242_141) begin
        banks_5_io_write_addr = _zz_io_write_addr_17;
      end
    end
    if(io_writeEn_18) begin
      if(when_BankedScratchMemory_l242_149) begin
        banks_5_io_write_addr = _zz_io_write_addr_18;
      end
    end
    if(io_writeEn_19) begin
      if(when_BankedScratchMemory_l242_157) begin
        banks_5_io_write_addr = _zz_io_write_addr_19;
      end
    end
    if(io_writeEn_20) begin
      if(when_BankedScratchMemory_l242_165) begin
        banks_5_io_write_addr = _zz_io_write_addr_20;
      end
    end
    if(io_writeEn_21) begin
      if(when_BankedScratchMemory_l242_173) begin
        banks_5_io_write_addr = _zz_io_write_addr_21;
      end
    end
    if(io_writeEn_22) begin
      if(when_BankedScratchMemory_l242_181) begin
        banks_5_io_write_addr = _zz_io_write_addr_22;
      end
    end
    if(io_writeEn_23) begin
      if(when_BankedScratchMemory_l242_189) begin
        banks_5_io_write_addr = _zz_io_write_addr_23;
      end
    end
    if(io_writeEn_24) begin
      if(when_BankedScratchMemory_l242_197) begin
        banks_5_io_write_addr = _zz_io_write_addr_24;
      end
    end
    if(io_writeEn_25) begin
      if(when_BankedScratchMemory_l242_205) begin
        banks_5_io_write_addr = _zz_io_write_addr_25;
      end
    end
    if(io_writeEn_26) begin
      if(when_BankedScratchMemory_l242_213) begin
        banks_5_io_write_addr = _zz_io_write_addr_26;
      end
    end
    if(io_writeEn_27) begin
      if(when_BankedScratchMemory_l242_221) begin
        banks_5_io_write_addr = _zz_io_write_addr_27;
      end
    end
  end

  always @(*) begin
    banks_5_io_write_data = 32'h0;
    if(io_writeEn_0) begin
      if(when_BankedScratchMemory_l242_5) begin
        banks_5_io_write_data = io_writeData_0;
      end
    end
    if(io_writeEn_1) begin
      if(when_BankedScratchMemory_l242_13) begin
        banks_5_io_write_data = io_writeData_1;
      end
    end
    if(io_writeEn_2) begin
      if(when_BankedScratchMemory_l242_21) begin
        banks_5_io_write_data = io_writeData_2;
      end
    end
    if(io_writeEn_3) begin
      if(when_BankedScratchMemory_l242_29) begin
        banks_5_io_write_data = io_writeData_3;
      end
    end
    if(io_writeEn_4) begin
      if(when_BankedScratchMemory_l242_37) begin
        banks_5_io_write_data = io_writeData_4;
      end
    end
    if(io_writeEn_5) begin
      if(when_BankedScratchMemory_l242_45) begin
        banks_5_io_write_data = io_writeData_5;
      end
    end
    if(io_writeEn_6) begin
      if(when_BankedScratchMemory_l242_53) begin
        banks_5_io_write_data = io_writeData_6;
      end
    end
    if(io_writeEn_7) begin
      if(when_BankedScratchMemory_l242_61) begin
        banks_5_io_write_data = io_writeData_7;
      end
    end
    if(io_writeEn_8) begin
      if(when_BankedScratchMemory_l242_69) begin
        banks_5_io_write_data = io_writeData_8;
      end
    end
    if(io_writeEn_9) begin
      if(when_BankedScratchMemory_l242_77) begin
        banks_5_io_write_data = io_writeData_9;
      end
    end
    if(io_writeEn_10) begin
      if(when_BankedScratchMemory_l242_85) begin
        banks_5_io_write_data = io_writeData_10;
      end
    end
    if(io_writeEn_11) begin
      if(when_BankedScratchMemory_l242_93) begin
        banks_5_io_write_data = io_writeData_11;
      end
    end
    if(io_writeEn_12) begin
      if(when_BankedScratchMemory_l242_101) begin
        banks_5_io_write_data = io_writeData_12;
      end
    end
    if(io_writeEn_13) begin
      if(when_BankedScratchMemory_l242_109) begin
        banks_5_io_write_data = io_writeData_13;
      end
    end
    if(io_writeEn_14) begin
      if(when_BankedScratchMemory_l242_117) begin
        banks_5_io_write_data = io_writeData_14;
      end
    end
    if(io_writeEn_15) begin
      if(when_BankedScratchMemory_l242_125) begin
        banks_5_io_write_data = io_writeData_15;
      end
    end
    if(io_writeEn_16) begin
      if(when_BankedScratchMemory_l242_133) begin
        banks_5_io_write_data = io_writeData_16;
      end
    end
    if(io_writeEn_17) begin
      if(when_BankedScratchMemory_l242_141) begin
        banks_5_io_write_data = io_writeData_17;
      end
    end
    if(io_writeEn_18) begin
      if(when_BankedScratchMemory_l242_149) begin
        banks_5_io_write_data = io_writeData_18;
      end
    end
    if(io_writeEn_19) begin
      if(when_BankedScratchMemory_l242_157) begin
        banks_5_io_write_data = io_writeData_19;
      end
    end
    if(io_writeEn_20) begin
      if(when_BankedScratchMemory_l242_165) begin
        banks_5_io_write_data = io_writeData_20;
      end
    end
    if(io_writeEn_21) begin
      if(when_BankedScratchMemory_l242_173) begin
        banks_5_io_write_data = io_writeData_21;
      end
    end
    if(io_writeEn_22) begin
      if(when_BankedScratchMemory_l242_181) begin
        banks_5_io_write_data = io_writeData_22;
      end
    end
    if(io_writeEn_23) begin
      if(when_BankedScratchMemory_l242_189) begin
        banks_5_io_write_data = io_writeData_23;
      end
    end
    if(io_writeEn_24) begin
      if(when_BankedScratchMemory_l242_197) begin
        banks_5_io_write_data = io_writeData_24;
      end
    end
    if(io_writeEn_25) begin
      if(when_BankedScratchMemory_l242_205) begin
        banks_5_io_write_data = io_writeData_25;
      end
    end
    if(io_writeEn_26) begin
      if(when_BankedScratchMemory_l242_213) begin
        banks_5_io_write_data = io_writeData_26;
      end
    end
    if(io_writeEn_27) begin
      if(when_BankedScratchMemory_l242_221) begin
        banks_5_io_write_data = io_writeData_27;
      end
    end
  end

  always @(*) begin
    banks_6_io_write_en = 1'b0;
    if(io_writeEn_0) begin
      if(when_BankedScratchMemory_l242_6) begin
        banks_6_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_1) begin
      if(when_BankedScratchMemory_l242_14) begin
        banks_6_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_2) begin
      if(when_BankedScratchMemory_l242_22) begin
        banks_6_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_3) begin
      if(when_BankedScratchMemory_l242_30) begin
        banks_6_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_4) begin
      if(when_BankedScratchMemory_l242_38) begin
        banks_6_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_5) begin
      if(when_BankedScratchMemory_l242_46) begin
        banks_6_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_6) begin
      if(when_BankedScratchMemory_l242_54) begin
        banks_6_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_7) begin
      if(when_BankedScratchMemory_l242_62) begin
        banks_6_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_8) begin
      if(when_BankedScratchMemory_l242_70) begin
        banks_6_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_9) begin
      if(when_BankedScratchMemory_l242_78) begin
        banks_6_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_10) begin
      if(when_BankedScratchMemory_l242_86) begin
        banks_6_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_11) begin
      if(when_BankedScratchMemory_l242_94) begin
        banks_6_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_12) begin
      if(when_BankedScratchMemory_l242_102) begin
        banks_6_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_13) begin
      if(when_BankedScratchMemory_l242_110) begin
        banks_6_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_14) begin
      if(when_BankedScratchMemory_l242_118) begin
        banks_6_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_15) begin
      if(when_BankedScratchMemory_l242_126) begin
        banks_6_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_16) begin
      if(when_BankedScratchMemory_l242_134) begin
        banks_6_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_17) begin
      if(when_BankedScratchMemory_l242_142) begin
        banks_6_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_18) begin
      if(when_BankedScratchMemory_l242_150) begin
        banks_6_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_19) begin
      if(when_BankedScratchMemory_l242_158) begin
        banks_6_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_20) begin
      if(when_BankedScratchMemory_l242_166) begin
        banks_6_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_21) begin
      if(when_BankedScratchMemory_l242_174) begin
        banks_6_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_22) begin
      if(when_BankedScratchMemory_l242_182) begin
        banks_6_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_23) begin
      if(when_BankedScratchMemory_l242_190) begin
        banks_6_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_24) begin
      if(when_BankedScratchMemory_l242_198) begin
        banks_6_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_25) begin
      if(when_BankedScratchMemory_l242_206) begin
        banks_6_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_26) begin
      if(when_BankedScratchMemory_l242_214) begin
        banks_6_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_27) begin
      if(when_BankedScratchMemory_l242_222) begin
        banks_6_io_write_en = 1'b1;
      end
    end
  end

  always @(*) begin
    banks_6_io_write_addr = 8'h0;
    if(io_writeEn_0) begin
      if(when_BankedScratchMemory_l242_6) begin
        banks_6_io_write_addr = _zz_io_write_addr;
      end
    end
    if(io_writeEn_1) begin
      if(when_BankedScratchMemory_l242_14) begin
        banks_6_io_write_addr = _zz_io_write_addr_1;
      end
    end
    if(io_writeEn_2) begin
      if(when_BankedScratchMemory_l242_22) begin
        banks_6_io_write_addr = _zz_io_write_addr_2;
      end
    end
    if(io_writeEn_3) begin
      if(when_BankedScratchMemory_l242_30) begin
        banks_6_io_write_addr = _zz_io_write_addr_3;
      end
    end
    if(io_writeEn_4) begin
      if(when_BankedScratchMemory_l242_38) begin
        banks_6_io_write_addr = _zz_io_write_addr_4;
      end
    end
    if(io_writeEn_5) begin
      if(when_BankedScratchMemory_l242_46) begin
        banks_6_io_write_addr = _zz_io_write_addr_5;
      end
    end
    if(io_writeEn_6) begin
      if(when_BankedScratchMemory_l242_54) begin
        banks_6_io_write_addr = _zz_io_write_addr_6;
      end
    end
    if(io_writeEn_7) begin
      if(when_BankedScratchMemory_l242_62) begin
        banks_6_io_write_addr = _zz_io_write_addr_7;
      end
    end
    if(io_writeEn_8) begin
      if(when_BankedScratchMemory_l242_70) begin
        banks_6_io_write_addr = _zz_io_write_addr_8;
      end
    end
    if(io_writeEn_9) begin
      if(when_BankedScratchMemory_l242_78) begin
        banks_6_io_write_addr = _zz_io_write_addr_9;
      end
    end
    if(io_writeEn_10) begin
      if(when_BankedScratchMemory_l242_86) begin
        banks_6_io_write_addr = _zz_io_write_addr_10;
      end
    end
    if(io_writeEn_11) begin
      if(when_BankedScratchMemory_l242_94) begin
        banks_6_io_write_addr = _zz_io_write_addr_11;
      end
    end
    if(io_writeEn_12) begin
      if(when_BankedScratchMemory_l242_102) begin
        banks_6_io_write_addr = _zz_io_write_addr_12;
      end
    end
    if(io_writeEn_13) begin
      if(when_BankedScratchMemory_l242_110) begin
        banks_6_io_write_addr = _zz_io_write_addr_13;
      end
    end
    if(io_writeEn_14) begin
      if(when_BankedScratchMemory_l242_118) begin
        banks_6_io_write_addr = _zz_io_write_addr_14;
      end
    end
    if(io_writeEn_15) begin
      if(when_BankedScratchMemory_l242_126) begin
        banks_6_io_write_addr = _zz_io_write_addr_15;
      end
    end
    if(io_writeEn_16) begin
      if(when_BankedScratchMemory_l242_134) begin
        banks_6_io_write_addr = _zz_io_write_addr_16;
      end
    end
    if(io_writeEn_17) begin
      if(when_BankedScratchMemory_l242_142) begin
        banks_6_io_write_addr = _zz_io_write_addr_17;
      end
    end
    if(io_writeEn_18) begin
      if(when_BankedScratchMemory_l242_150) begin
        banks_6_io_write_addr = _zz_io_write_addr_18;
      end
    end
    if(io_writeEn_19) begin
      if(when_BankedScratchMemory_l242_158) begin
        banks_6_io_write_addr = _zz_io_write_addr_19;
      end
    end
    if(io_writeEn_20) begin
      if(when_BankedScratchMemory_l242_166) begin
        banks_6_io_write_addr = _zz_io_write_addr_20;
      end
    end
    if(io_writeEn_21) begin
      if(when_BankedScratchMemory_l242_174) begin
        banks_6_io_write_addr = _zz_io_write_addr_21;
      end
    end
    if(io_writeEn_22) begin
      if(when_BankedScratchMemory_l242_182) begin
        banks_6_io_write_addr = _zz_io_write_addr_22;
      end
    end
    if(io_writeEn_23) begin
      if(when_BankedScratchMemory_l242_190) begin
        banks_6_io_write_addr = _zz_io_write_addr_23;
      end
    end
    if(io_writeEn_24) begin
      if(when_BankedScratchMemory_l242_198) begin
        banks_6_io_write_addr = _zz_io_write_addr_24;
      end
    end
    if(io_writeEn_25) begin
      if(when_BankedScratchMemory_l242_206) begin
        banks_6_io_write_addr = _zz_io_write_addr_25;
      end
    end
    if(io_writeEn_26) begin
      if(when_BankedScratchMemory_l242_214) begin
        banks_6_io_write_addr = _zz_io_write_addr_26;
      end
    end
    if(io_writeEn_27) begin
      if(when_BankedScratchMemory_l242_222) begin
        banks_6_io_write_addr = _zz_io_write_addr_27;
      end
    end
  end

  always @(*) begin
    banks_6_io_write_data = 32'h0;
    if(io_writeEn_0) begin
      if(when_BankedScratchMemory_l242_6) begin
        banks_6_io_write_data = io_writeData_0;
      end
    end
    if(io_writeEn_1) begin
      if(when_BankedScratchMemory_l242_14) begin
        banks_6_io_write_data = io_writeData_1;
      end
    end
    if(io_writeEn_2) begin
      if(when_BankedScratchMemory_l242_22) begin
        banks_6_io_write_data = io_writeData_2;
      end
    end
    if(io_writeEn_3) begin
      if(when_BankedScratchMemory_l242_30) begin
        banks_6_io_write_data = io_writeData_3;
      end
    end
    if(io_writeEn_4) begin
      if(when_BankedScratchMemory_l242_38) begin
        banks_6_io_write_data = io_writeData_4;
      end
    end
    if(io_writeEn_5) begin
      if(when_BankedScratchMemory_l242_46) begin
        banks_6_io_write_data = io_writeData_5;
      end
    end
    if(io_writeEn_6) begin
      if(when_BankedScratchMemory_l242_54) begin
        banks_6_io_write_data = io_writeData_6;
      end
    end
    if(io_writeEn_7) begin
      if(when_BankedScratchMemory_l242_62) begin
        banks_6_io_write_data = io_writeData_7;
      end
    end
    if(io_writeEn_8) begin
      if(when_BankedScratchMemory_l242_70) begin
        banks_6_io_write_data = io_writeData_8;
      end
    end
    if(io_writeEn_9) begin
      if(when_BankedScratchMemory_l242_78) begin
        banks_6_io_write_data = io_writeData_9;
      end
    end
    if(io_writeEn_10) begin
      if(when_BankedScratchMemory_l242_86) begin
        banks_6_io_write_data = io_writeData_10;
      end
    end
    if(io_writeEn_11) begin
      if(when_BankedScratchMemory_l242_94) begin
        banks_6_io_write_data = io_writeData_11;
      end
    end
    if(io_writeEn_12) begin
      if(when_BankedScratchMemory_l242_102) begin
        banks_6_io_write_data = io_writeData_12;
      end
    end
    if(io_writeEn_13) begin
      if(when_BankedScratchMemory_l242_110) begin
        banks_6_io_write_data = io_writeData_13;
      end
    end
    if(io_writeEn_14) begin
      if(when_BankedScratchMemory_l242_118) begin
        banks_6_io_write_data = io_writeData_14;
      end
    end
    if(io_writeEn_15) begin
      if(when_BankedScratchMemory_l242_126) begin
        banks_6_io_write_data = io_writeData_15;
      end
    end
    if(io_writeEn_16) begin
      if(when_BankedScratchMemory_l242_134) begin
        banks_6_io_write_data = io_writeData_16;
      end
    end
    if(io_writeEn_17) begin
      if(when_BankedScratchMemory_l242_142) begin
        banks_6_io_write_data = io_writeData_17;
      end
    end
    if(io_writeEn_18) begin
      if(when_BankedScratchMemory_l242_150) begin
        banks_6_io_write_data = io_writeData_18;
      end
    end
    if(io_writeEn_19) begin
      if(when_BankedScratchMemory_l242_158) begin
        banks_6_io_write_data = io_writeData_19;
      end
    end
    if(io_writeEn_20) begin
      if(when_BankedScratchMemory_l242_166) begin
        banks_6_io_write_data = io_writeData_20;
      end
    end
    if(io_writeEn_21) begin
      if(when_BankedScratchMemory_l242_174) begin
        banks_6_io_write_data = io_writeData_21;
      end
    end
    if(io_writeEn_22) begin
      if(when_BankedScratchMemory_l242_182) begin
        banks_6_io_write_data = io_writeData_22;
      end
    end
    if(io_writeEn_23) begin
      if(when_BankedScratchMemory_l242_190) begin
        banks_6_io_write_data = io_writeData_23;
      end
    end
    if(io_writeEn_24) begin
      if(when_BankedScratchMemory_l242_198) begin
        banks_6_io_write_data = io_writeData_24;
      end
    end
    if(io_writeEn_25) begin
      if(when_BankedScratchMemory_l242_206) begin
        banks_6_io_write_data = io_writeData_25;
      end
    end
    if(io_writeEn_26) begin
      if(when_BankedScratchMemory_l242_214) begin
        banks_6_io_write_data = io_writeData_26;
      end
    end
    if(io_writeEn_27) begin
      if(when_BankedScratchMemory_l242_222) begin
        banks_6_io_write_data = io_writeData_27;
      end
    end
  end

  always @(*) begin
    banks_7_io_write_en = 1'b0;
    if(io_writeEn_0) begin
      if(when_BankedScratchMemory_l242_7) begin
        banks_7_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_1) begin
      if(when_BankedScratchMemory_l242_15) begin
        banks_7_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_2) begin
      if(when_BankedScratchMemory_l242_23) begin
        banks_7_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_3) begin
      if(when_BankedScratchMemory_l242_31) begin
        banks_7_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_4) begin
      if(when_BankedScratchMemory_l242_39) begin
        banks_7_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_5) begin
      if(when_BankedScratchMemory_l242_47) begin
        banks_7_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_6) begin
      if(when_BankedScratchMemory_l242_55) begin
        banks_7_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_7) begin
      if(when_BankedScratchMemory_l242_63) begin
        banks_7_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_8) begin
      if(when_BankedScratchMemory_l242_71) begin
        banks_7_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_9) begin
      if(when_BankedScratchMemory_l242_79) begin
        banks_7_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_10) begin
      if(when_BankedScratchMemory_l242_87) begin
        banks_7_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_11) begin
      if(when_BankedScratchMemory_l242_95) begin
        banks_7_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_12) begin
      if(when_BankedScratchMemory_l242_103) begin
        banks_7_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_13) begin
      if(when_BankedScratchMemory_l242_111) begin
        banks_7_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_14) begin
      if(when_BankedScratchMemory_l242_119) begin
        banks_7_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_15) begin
      if(when_BankedScratchMemory_l242_127) begin
        banks_7_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_16) begin
      if(when_BankedScratchMemory_l242_135) begin
        banks_7_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_17) begin
      if(when_BankedScratchMemory_l242_143) begin
        banks_7_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_18) begin
      if(when_BankedScratchMemory_l242_151) begin
        banks_7_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_19) begin
      if(when_BankedScratchMemory_l242_159) begin
        banks_7_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_20) begin
      if(when_BankedScratchMemory_l242_167) begin
        banks_7_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_21) begin
      if(when_BankedScratchMemory_l242_175) begin
        banks_7_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_22) begin
      if(when_BankedScratchMemory_l242_183) begin
        banks_7_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_23) begin
      if(when_BankedScratchMemory_l242_191) begin
        banks_7_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_24) begin
      if(when_BankedScratchMemory_l242_199) begin
        banks_7_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_25) begin
      if(when_BankedScratchMemory_l242_207) begin
        banks_7_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_26) begin
      if(when_BankedScratchMemory_l242_215) begin
        banks_7_io_write_en = 1'b1;
      end
    end
    if(io_writeEn_27) begin
      if(when_BankedScratchMemory_l242_223) begin
        banks_7_io_write_en = 1'b1;
      end
    end
  end

  always @(*) begin
    banks_7_io_write_addr = 8'h0;
    if(io_writeEn_0) begin
      if(when_BankedScratchMemory_l242_7) begin
        banks_7_io_write_addr = _zz_io_write_addr;
      end
    end
    if(io_writeEn_1) begin
      if(when_BankedScratchMemory_l242_15) begin
        banks_7_io_write_addr = _zz_io_write_addr_1;
      end
    end
    if(io_writeEn_2) begin
      if(when_BankedScratchMemory_l242_23) begin
        banks_7_io_write_addr = _zz_io_write_addr_2;
      end
    end
    if(io_writeEn_3) begin
      if(when_BankedScratchMemory_l242_31) begin
        banks_7_io_write_addr = _zz_io_write_addr_3;
      end
    end
    if(io_writeEn_4) begin
      if(when_BankedScratchMemory_l242_39) begin
        banks_7_io_write_addr = _zz_io_write_addr_4;
      end
    end
    if(io_writeEn_5) begin
      if(when_BankedScratchMemory_l242_47) begin
        banks_7_io_write_addr = _zz_io_write_addr_5;
      end
    end
    if(io_writeEn_6) begin
      if(when_BankedScratchMemory_l242_55) begin
        banks_7_io_write_addr = _zz_io_write_addr_6;
      end
    end
    if(io_writeEn_7) begin
      if(when_BankedScratchMemory_l242_63) begin
        banks_7_io_write_addr = _zz_io_write_addr_7;
      end
    end
    if(io_writeEn_8) begin
      if(when_BankedScratchMemory_l242_71) begin
        banks_7_io_write_addr = _zz_io_write_addr_8;
      end
    end
    if(io_writeEn_9) begin
      if(when_BankedScratchMemory_l242_79) begin
        banks_7_io_write_addr = _zz_io_write_addr_9;
      end
    end
    if(io_writeEn_10) begin
      if(when_BankedScratchMemory_l242_87) begin
        banks_7_io_write_addr = _zz_io_write_addr_10;
      end
    end
    if(io_writeEn_11) begin
      if(when_BankedScratchMemory_l242_95) begin
        banks_7_io_write_addr = _zz_io_write_addr_11;
      end
    end
    if(io_writeEn_12) begin
      if(when_BankedScratchMemory_l242_103) begin
        banks_7_io_write_addr = _zz_io_write_addr_12;
      end
    end
    if(io_writeEn_13) begin
      if(when_BankedScratchMemory_l242_111) begin
        banks_7_io_write_addr = _zz_io_write_addr_13;
      end
    end
    if(io_writeEn_14) begin
      if(when_BankedScratchMemory_l242_119) begin
        banks_7_io_write_addr = _zz_io_write_addr_14;
      end
    end
    if(io_writeEn_15) begin
      if(when_BankedScratchMemory_l242_127) begin
        banks_7_io_write_addr = _zz_io_write_addr_15;
      end
    end
    if(io_writeEn_16) begin
      if(when_BankedScratchMemory_l242_135) begin
        banks_7_io_write_addr = _zz_io_write_addr_16;
      end
    end
    if(io_writeEn_17) begin
      if(when_BankedScratchMemory_l242_143) begin
        banks_7_io_write_addr = _zz_io_write_addr_17;
      end
    end
    if(io_writeEn_18) begin
      if(when_BankedScratchMemory_l242_151) begin
        banks_7_io_write_addr = _zz_io_write_addr_18;
      end
    end
    if(io_writeEn_19) begin
      if(when_BankedScratchMemory_l242_159) begin
        banks_7_io_write_addr = _zz_io_write_addr_19;
      end
    end
    if(io_writeEn_20) begin
      if(when_BankedScratchMemory_l242_167) begin
        banks_7_io_write_addr = _zz_io_write_addr_20;
      end
    end
    if(io_writeEn_21) begin
      if(when_BankedScratchMemory_l242_175) begin
        banks_7_io_write_addr = _zz_io_write_addr_21;
      end
    end
    if(io_writeEn_22) begin
      if(when_BankedScratchMemory_l242_183) begin
        banks_7_io_write_addr = _zz_io_write_addr_22;
      end
    end
    if(io_writeEn_23) begin
      if(when_BankedScratchMemory_l242_191) begin
        banks_7_io_write_addr = _zz_io_write_addr_23;
      end
    end
    if(io_writeEn_24) begin
      if(when_BankedScratchMemory_l242_199) begin
        banks_7_io_write_addr = _zz_io_write_addr_24;
      end
    end
    if(io_writeEn_25) begin
      if(when_BankedScratchMemory_l242_207) begin
        banks_7_io_write_addr = _zz_io_write_addr_25;
      end
    end
    if(io_writeEn_26) begin
      if(when_BankedScratchMemory_l242_215) begin
        banks_7_io_write_addr = _zz_io_write_addr_26;
      end
    end
    if(io_writeEn_27) begin
      if(when_BankedScratchMemory_l242_223) begin
        banks_7_io_write_addr = _zz_io_write_addr_27;
      end
    end
  end

  always @(*) begin
    banks_7_io_write_data = 32'h0;
    if(io_writeEn_0) begin
      if(when_BankedScratchMemory_l242_7) begin
        banks_7_io_write_data = io_writeData_0;
      end
    end
    if(io_writeEn_1) begin
      if(when_BankedScratchMemory_l242_15) begin
        banks_7_io_write_data = io_writeData_1;
      end
    end
    if(io_writeEn_2) begin
      if(when_BankedScratchMemory_l242_23) begin
        banks_7_io_write_data = io_writeData_2;
      end
    end
    if(io_writeEn_3) begin
      if(when_BankedScratchMemory_l242_31) begin
        banks_7_io_write_data = io_writeData_3;
      end
    end
    if(io_writeEn_4) begin
      if(when_BankedScratchMemory_l242_39) begin
        banks_7_io_write_data = io_writeData_4;
      end
    end
    if(io_writeEn_5) begin
      if(when_BankedScratchMemory_l242_47) begin
        banks_7_io_write_data = io_writeData_5;
      end
    end
    if(io_writeEn_6) begin
      if(when_BankedScratchMemory_l242_55) begin
        banks_7_io_write_data = io_writeData_6;
      end
    end
    if(io_writeEn_7) begin
      if(when_BankedScratchMemory_l242_63) begin
        banks_7_io_write_data = io_writeData_7;
      end
    end
    if(io_writeEn_8) begin
      if(when_BankedScratchMemory_l242_71) begin
        banks_7_io_write_data = io_writeData_8;
      end
    end
    if(io_writeEn_9) begin
      if(when_BankedScratchMemory_l242_79) begin
        banks_7_io_write_data = io_writeData_9;
      end
    end
    if(io_writeEn_10) begin
      if(when_BankedScratchMemory_l242_87) begin
        banks_7_io_write_data = io_writeData_10;
      end
    end
    if(io_writeEn_11) begin
      if(when_BankedScratchMemory_l242_95) begin
        banks_7_io_write_data = io_writeData_11;
      end
    end
    if(io_writeEn_12) begin
      if(when_BankedScratchMemory_l242_103) begin
        banks_7_io_write_data = io_writeData_12;
      end
    end
    if(io_writeEn_13) begin
      if(when_BankedScratchMemory_l242_111) begin
        banks_7_io_write_data = io_writeData_13;
      end
    end
    if(io_writeEn_14) begin
      if(when_BankedScratchMemory_l242_119) begin
        banks_7_io_write_data = io_writeData_14;
      end
    end
    if(io_writeEn_15) begin
      if(when_BankedScratchMemory_l242_127) begin
        banks_7_io_write_data = io_writeData_15;
      end
    end
    if(io_writeEn_16) begin
      if(when_BankedScratchMemory_l242_135) begin
        banks_7_io_write_data = io_writeData_16;
      end
    end
    if(io_writeEn_17) begin
      if(when_BankedScratchMemory_l242_143) begin
        banks_7_io_write_data = io_writeData_17;
      end
    end
    if(io_writeEn_18) begin
      if(when_BankedScratchMemory_l242_151) begin
        banks_7_io_write_data = io_writeData_18;
      end
    end
    if(io_writeEn_19) begin
      if(when_BankedScratchMemory_l242_159) begin
        banks_7_io_write_data = io_writeData_19;
      end
    end
    if(io_writeEn_20) begin
      if(when_BankedScratchMemory_l242_167) begin
        banks_7_io_write_data = io_writeData_20;
      end
    end
    if(io_writeEn_21) begin
      if(when_BankedScratchMemory_l242_175) begin
        banks_7_io_write_data = io_writeData_21;
      end
    end
    if(io_writeEn_22) begin
      if(when_BankedScratchMemory_l242_183) begin
        banks_7_io_write_data = io_writeData_22;
      end
    end
    if(io_writeEn_23) begin
      if(when_BankedScratchMemory_l242_191) begin
        banks_7_io_write_data = io_writeData_23;
      end
    end
    if(io_writeEn_24) begin
      if(when_BankedScratchMemory_l242_199) begin
        banks_7_io_write_data = io_writeData_24;
      end
    end
    if(io_writeEn_25) begin
      if(when_BankedScratchMemory_l242_207) begin
        banks_7_io_write_data = io_writeData_25;
      end
    end
    if(io_writeEn_26) begin
      if(when_BankedScratchMemory_l242_215) begin
        banks_7_io_write_data = io_writeData_26;
      end
    end
    if(io_writeEn_27) begin
      if(when_BankedScratchMemory_l242_223) begin
        banks_7_io_write_data = io_writeData_27;
      end
    end
  end

  assign _zz_when_BankedScratchMemory_l242 = io_writeAddr_0[2 : 0];
  assign _zz_io_write_addr = io_writeAddr_0[10 : 3];
  assign when_BankedScratchMemory_l242 = (_zz_when_BankedScratchMemory_l242 == 3'b000);
  assign when_BankedScratchMemory_l242_1 = (_zz_when_BankedScratchMemory_l242 == 3'b001);
  assign when_BankedScratchMemory_l242_2 = (_zz_when_BankedScratchMemory_l242 == 3'b010);
  assign when_BankedScratchMemory_l242_3 = (_zz_when_BankedScratchMemory_l242 == 3'b011);
  assign when_BankedScratchMemory_l242_4 = (_zz_when_BankedScratchMemory_l242 == 3'b100);
  assign when_BankedScratchMemory_l242_5 = (_zz_when_BankedScratchMemory_l242 == 3'b101);
  assign when_BankedScratchMemory_l242_6 = (_zz_when_BankedScratchMemory_l242 == 3'b110);
  assign when_BankedScratchMemory_l242_7 = (_zz_when_BankedScratchMemory_l242 == 3'b111);
  assign _zz_when_BankedScratchMemory_l242_1 = io_writeAddr_1[2 : 0];
  assign _zz_io_write_addr_1 = io_writeAddr_1[10 : 3];
  assign when_BankedScratchMemory_l242_8 = (_zz_when_BankedScratchMemory_l242_1 == 3'b000);
  assign when_BankedScratchMemory_l242_9 = (_zz_when_BankedScratchMemory_l242_1 == 3'b001);
  assign when_BankedScratchMemory_l242_10 = (_zz_when_BankedScratchMemory_l242_1 == 3'b010);
  assign when_BankedScratchMemory_l242_11 = (_zz_when_BankedScratchMemory_l242_1 == 3'b011);
  assign when_BankedScratchMemory_l242_12 = (_zz_when_BankedScratchMemory_l242_1 == 3'b100);
  assign when_BankedScratchMemory_l242_13 = (_zz_when_BankedScratchMemory_l242_1 == 3'b101);
  assign when_BankedScratchMemory_l242_14 = (_zz_when_BankedScratchMemory_l242_1 == 3'b110);
  assign when_BankedScratchMemory_l242_15 = (_zz_when_BankedScratchMemory_l242_1 == 3'b111);
  assign _zz_when_BankedScratchMemory_l242_2 = io_writeAddr_2[2 : 0];
  assign _zz_io_write_addr_2 = io_writeAddr_2[10 : 3];
  assign when_BankedScratchMemory_l242_16 = (_zz_when_BankedScratchMemory_l242_2 == 3'b000);
  assign when_BankedScratchMemory_l242_17 = (_zz_when_BankedScratchMemory_l242_2 == 3'b001);
  assign when_BankedScratchMemory_l242_18 = (_zz_when_BankedScratchMemory_l242_2 == 3'b010);
  assign when_BankedScratchMemory_l242_19 = (_zz_when_BankedScratchMemory_l242_2 == 3'b011);
  assign when_BankedScratchMemory_l242_20 = (_zz_when_BankedScratchMemory_l242_2 == 3'b100);
  assign when_BankedScratchMemory_l242_21 = (_zz_when_BankedScratchMemory_l242_2 == 3'b101);
  assign when_BankedScratchMemory_l242_22 = (_zz_when_BankedScratchMemory_l242_2 == 3'b110);
  assign when_BankedScratchMemory_l242_23 = (_zz_when_BankedScratchMemory_l242_2 == 3'b111);
  assign _zz_when_BankedScratchMemory_l242_3 = io_writeAddr_3[2 : 0];
  assign _zz_io_write_addr_3 = io_writeAddr_3[10 : 3];
  assign when_BankedScratchMemory_l242_24 = (_zz_when_BankedScratchMemory_l242_3 == 3'b000);
  assign when_BankedScratchMemory_l242_25 = (_zz_when_BankedScratchMemory_l242_3 == 3'b001);
  assign when_BankedScratchMemory_l242_26 = (_zz_when_BankedScratchMemory_l242_3 == 3'b010);
  assign when_BankedScratchMemory_l242_27 = (_zz_when_BankedScratchMemory_l242_3 == 3'b011);
  assign when_BankedScratchMemory_l242_28 = (_zz_when_BankedScratchMemory_l242_3 == 3'b100);
  assign when_BankedScratchMemory_l242_29 = (_zz_when_BankedScratchMemory_l242_3 == 3'b101);
  assign when_BankedScratchMemory_l242_30 = (_zz_when_BankedScratchMemory_l242_3 == 3'b110);
  assign when_BankedScratchMemory_l242_31 = (_zz_when_BankedScratchMemory_l242_3 == 3'b111);
  assign _zz_when_BankedScratchMemory_l242_4 = io_writeAddr_4[2 : 0];
  assign _zz_io_write_addr_4 = io_writeAddr_4[10 : 3];
  assign when_BankedScratchMemory_l242_32 = (_zz_when_BankedScratchMemory_l242_4 == 3'b000);
  assign when_BankedScratchMemory_l242_33 = (_zz_when_BankedScratchMemory_l242_4 == 3'b001);
  assign when_BankedScratchMemory_l242_34 = (_zz_when_BankedScratchMemory_l242_4 == 3'b010);
  assign when_BankedScratchMemory_l242_35 = (_zz_when_BankedScratchMemory_l242_4 == 3'b011);
  assign when_BankedScratchMemory_l242_36 = (_zz_when_BankedScratchMemory_l242_4 == 3'b100);
  assign when_BankedScratchMemory_l242_37 = (_zz_when_BankedScratchMemory_l242_4 == 3'b101);
  assign when_BankedScratchMemory_l242_38 = (_zz_when_BankedScratchMemory_l242_4 == 3'b110);
  assign when_BankedScratchMemory_l242_39 = (_zz_when_BankedScratchMemory_l242_4 == 3'b111);
  assign _zz_when_BankedScratchMemory_l242_5 = io_writeAddr_5[2 : 0];
  assign _zz_io_write_addr_5 = io_writeAddr_5[10 : 3];
  assign when_BankedScratchMemory_l242_40 = (_zz_when_BankedScratchMemory_l242_5 == 3'b000);
  assign when_BankedScratchMemory_l242_41 = (_zz_when_BankedScratchMemory_l242_5 == 3'b001);
  assign when_BankedScratchMemory_l242_42 = (_zz_when_BankedScratchMemory_l242_5 == 3'b010);
  assign when_BankedScratchMemory_l242_43 = (_zz_when_BankedScratchMemory_l242_5 == 3'b011);
  assign when_BankedScratchMemory_l242_44 = (_zz_when_BankedScratchMemory_l242_5 == 3'b100);
  assign when_BankedScratchMemory_l242_45 = (_zz_when_BankedScratchMemory_l242_5 == 3'b101);
  assign when_BankedScratchMemory_l242_46 = (_zz_when_BankedScratchMemory_l242_5 == 3'b110);
  assign when_BankedScratchMemory_l242_47 = (_zz_when_BankedScratchMemory_l242_5 == 3'b111);
  assign _zz_when_BankedScratchMemory_l242_6 = io_writeAddr_6[2 : 0];
  assign _zz_io_write_addr_6 = io_writeAddr_6[10 : 3];
  assign when_BankedScratchMemory_l242_48 = (_zz_when_BankedScratchMemory_l242_6 == 3'b000);
  assign when_BankedScratchMemory_l242_49 = (_zz_when_BankedScratchMemory_l242_6 == 3'b001);
  assign when_BankedScratchMemory_l242_50 = (_zz_when_BankedScratchMemory_l242_6 == 3'b010);
  assign when_BankedScratchMemory_l242_51 = (_zz_when_BankedScratchMemory_l242_6 == 3'b011);
  assign when_BankedScratchMemory_l242_52 = (_zz_when_BankedScratchMemory_l242_6 == 3'b100);
  assign when_BankedScratchMemory_l242_53 = (_zz_when_BankedScratchMemory_l242_6 == 3'b101);
  assign when_BankedScratchMemory_l242_54 = (_zz_when_BankedScratchMemory_l242_6 == 3'b110);
  assign when_BankedScratchMemory_l242_55 = (_zz_when_BankedScratchMemory_l242_6 == 3'b111);
  assign _zz_when_BankedScratchMemory_l242_7 = io_writeAddr_7[2 : 0];
  assign _zz_io_write_addr_7 = io_writeAddr_7[10 : 3];
  assign when_BankedScratchMemory_l242_56 = (_zz_when_BankedScratchMemory_l242_7 == 3'b000);
  assign when_BankedScratchMemory_l242_57 = (_zz_when_BankedScratchMemory_l242_7 == 3'b001);
  assign when_BankedScratchMemory_l242_58 = (_zz_when_BankedScratchMemory_l242_7 == 3'b010);
  assign when_BankedScratchMemory_l242_59 = (_zz_when_BankedScratchMemory_l242_7 == 3'b011);
  assign when_BankedScratchMemory_l242_60 = (_zz_when_BankedScratchMemory_l242_7 == 3'b100);
  assign when_BankedScratchMemory_l242_61 = (_zz_when_BankedScratchMemory_l242_7 == 3'b101);
  assign when_BankedScratchMemory_l242_62 = (_zz_when_BankedScratchMemory_l242_7 == 3'b110);
  assign when_BankedScratchMemory_l242_63 = (_zz_when_BankedScratchMemory_l242_7 == 3'b111);
  assign _zz_when_BankedScratchMemory_l242_8 = io_writeAddr_8[2 : 0];
  assign _zz_io_write_addr_8 = io_writeAddr_8[10 : 3];
  assign when_BankedScratchMemory_l242_64 = (_zz_when_BankedScratchMemory_l242_8 == 3'b000);
  assign when_BankedScratchMemory_l242_65 = (_zz_when_BankedScratchMemory_l242_8 == 3'b001);
  assign when_BankedScratchMemory_l242_66 = (_zz_when_BankedScratchMemory_l242_8 == 3'b010);
  assign when_BankedScratchMemory_l242_67 = (_zz_when_BankedScratchMemory_l242_8 == 3'b011);
  assign when_BankedScratchMemory_l242_68 = (_zz_when_BankedScratchMemory_l242_8 == 3'b100);
  assign when_BankedScratchMemory_l242_69 = (_zz_when_BankedScratchMemory_l242_8 == 3'b101);
  assign when_BankedScratchMemory_l242_70 = (_zz_when_BankedScratchMemory_l242_8 == 3'b110);
  assign when_BankedScratchMemory_l242_71 = (_zz_when_BankedScratchMemory_l242_8 == 3'b111);
  assign _zz_when_BankedScratchMemory_l242_9 = io_writeAddr_9[2 : 0];
  assign _zz_io_write_addr_9 = io_writeAddr_9[10 : 3];
  assign when_BankedScratchMemory_l242_72 = (_zz_when_BankedScratchMemory_l242_9 == 3'b000);
  assign when_BankedScratchMemory_l242_73 = (_zz_when_BankedScratchMemory_l242_9 == 3'b001);
  assign when_BankedScratchMemory_l242_74 = (_zz_when_BankedScratchMemory_l242_9 == 3'b010);
  assign when_BankedScratchMemory_l242_75 = (_zz_when_BankedScratchMemory_l242_9 == 3'b011);
  assign when_BankedScratchMemory_l242_76 = (_zz_when_BankedScratchMemory_l242_9 == 3'b100);
  assign when_BankedScratchMemory_l242_77 = (_zz_when_BankedScratchMemory_l242_9 == 3'b101);
  assign when_BankedScratchMemory_l242_78 = (_zz_when_BankedScratchMemory_l242_9 == 3'b110);
  assign when_BankedScratchMemory_l242_79 = (_zz_when_BankedScratchMemory_l242_9 == 3'b111);
  assign _zz_when_BankedScratchMemory_l242_10 = io_writeAddr_10[2 : 0];
  assign _zz_io_write_addr_10 = io_writeAddr_10[10 : 3];
  assign when_BankedScratchMemory_l242_80 = (_zz_when_BankedScratchMemory_l242_10 == 3'b000);
  assign when_BankedScratchMemory_l242_81 = (_zz_when_BankedScratchMemory_l242_10 == 3'b001);
  assign when_BankedScratchMemory_l242_82 = (_zz_when_BankedScratchMemory_l242_10 == 3'b010);
  assign when_BankedScratchMemory_l242_83 = (_zz_when_BankedScratchMemory_l242_10 == 3'b011);
  assign when_BankedScratchMemory_l242_84 = (_zz_when_BankedScratchMemory_l242_10 == 3'b100);
  assign when_BankedScratchMemory_l242_85 = (_zz_when_BankedScratchMemory_l242_10 == 3'b101);
  assign when_BankedScratchMemory_l242_86 = (_zz_when_BankedScratchMemory_l242_10 == 3'b110);
  assign when_BankedScratchMemory_l242_87 = (_zz_when_BankedScratchMemory_l242_10 == 3'b111);
  assign _zz_when_BankedScratchMemory_l242_11 = io_writeAddr_11[2 : 0];
  assign _zz_io_write_addr_11 = io_writeAddr_11[10 : 3];
  assign when_BankedScratchMemory_l242_88 = (_zz_when_BankedScratchMemory_l242_11 == 3'b000);
  assign when_BankedScratchMemory_l242_89 = (_zz_when_BankedScratchMemory_l242_11 == 3'b001);
  assign when_BankedScratchMemory_l242_90 = (_zz_when_BankedScratchMemory_l242_11 == 3'b010);
  assign when_BankedScratchMemory_l242_91 = (_zz_when_BankedScratchMemory_l242_11 == 3'b011);
  assign when_BankedScratchMemory_l242_92 = (_zz_when_BankedScratchMemory_l242_11 == 3'b100);
  assign when_BankedScratchMemory_l242_93 = (_zz_when_BankedScratchMemory_l242_11 == 3'b101);
  assign when_BankedScratchMemory_l242_94 = (_zz_when_BankedScratchMemory_l242_11 == 3'b110);
  assign when_BankedScratchMemory_l242_95 = (_zz_when_BankedScratchMemory_l242_11 == 3'b111);
  assign _zz_when_BankedScratchMemory_l242_12 = io_writeAddr_12[2 : 0];
  assign _zz_io_write_addr_12 = io_writeAddr_12[10 : 3];
  assign when_BankedScratchMemory_l242_96 = (_zz_when_BankedScratchMemory_l242_12 == 3'b000);
  assign when_BankedScratchMemory_l242_97 = (_zz_when_BankedScratchMemory_l242_12 == 3'b001);
  assign when_BankedScratchMemory_l242_98 = (_zz_when_BankedScratchMemory_l242_12 == 3'b010);
  assign when_BankedScratchMemory_l242_99 = (_zz_when_BankedScratchMemory_l242_12 == 3'b011);
  assign when_BankedScratchMemory_l242_100 = (_zz_when_BankedScratchMemory_l242_12 == 3'b100);
  assign when_BankedScratchMemory_l242_101 = (_zz_when_BankedScratchMemory_l242_12 == 3'b101);
  assign when_BankedScratchMemory_l242_102 = (_zz_when_BankedScratchMemory_l242_12 == 3'b110);
  assign when_BankedScratchMemory_l242_103 = (_zz_when_BankedScratchMemory_l242_12 == 3'b111);
  assign _zz_when_BankedScratchMemory_l242_13 = io_writeAddr_13[2 : 0];
  assign _zz_io_write_addr_13 = io_writeAddr_13[10 : 3];
  assign when_BankedScratchMemory_l242_104 = (_zz_when_BankedScratchMemory_l242_13 == 3'b000);
  assign when_BankedScratchMemory_l242_105 = (_zz_when_BankedScratchMemory_l242_13 == 3'b001);
  assign when_BankedScratchMemory_l242_106 = (_zz_when_BankedScratchMemory_l242_13 == 3'b010);
  assign when_BankedScratchMemory_l242_107 = (_zz_when_BankedScratchMemory_l242_13 == 3'b011);
  assign when_BankedScratchMemory_l242_108 = (_zz_when_BankedScratchMemory_l242_13 == 3'b100);
  assign when_BankedScratchMemory_l242_109 = (_zz_when_BankedScratchMemory_l242_13 == 3'b101);
  assign when_BankedScratchMemory_l242_110 = (_zz_when_BankedScratchMemory_l242_13 == 3'b110);
  assign when_BankedScratchMemory_l242_111 = (_zz_when_BankedScratchMemory_l242_13 == 3'b111);
  assign _zz_when_BankedScratchMemory_l242_14 = io_writeAddr_14[2 : 0];
  assign _zz_io_write_addr_14 = io_writeAddr_14[10 : 3];
  assign when_BankedScratchMemory_l242_112 = (_zz_when_BankedScratchMemory_l242_14 == 3'b000);
  assign when_BankedScratchMemory_l242_113 = (_zz_when_BankedScratchMemory_l242_14 == 3'b001);
  assign when_BankedScratchMemory_l242_114 = (_zz_when_BankedScratchMemory_l242_14 == 3'b010);
  assign when_BankedScratchMemory_l242_115 = (_zz_when_BankedScratchMemory_l242_14 == 3'b011);
  assign when_BankedScratchMemory_l242_116 = (_zz_when_BankedScratchMemory_l242_14 == 3'b100);
  assign when_BankedScratchMemory_l242_117 = (_zz_when_BankedScratchMemory_l242_14 == 3'b101);
  assign when_BankedScratchMemory_l242_118 = (_zz_when_BankedScratchMemory_l242_14 == 3'b110);
  assign when_BankedScratchMemory_l242_119 = (_zz_when_BankedScratchMemory_l242_14 == 3'b111);
  assign _zz_when_BankedScratchMemory_l242_15 = io_writeAddr_15[2 : 0];
  assign _zz_io_write_addr_15 = io_writeAddr_15[10 : 3];
  assign when_BankedScratchMemory_l242_120 = (_zz_when_BankedScratchMemory_l242_15 == 3'b000);
  assign when_BankedScratchMemory_l242_121 = (_zz_when_BankedScratchMemory_l242_15 == 3'b001);
  assign when_BankedScratchMemory_l242_122 = (_zz_when_BankedScratchMemory_l242_15 == 3'b010);
  assign when_BankedScratchMemory_l242_123 = (_zz_when_BankedScratchMemory_l242_15 == 3'b011);
  assign when_BankedScratchMemory_l242_124 = (_zz_when_BankedScratchMemory_l242_15 == 3'b100);
  assign when_BankedScratchMemory_l242_125 = (_zz_when_BankedScratchMemory_l242_15 == 3'b101);
  assign when_BankedScratchMemory_l242_126 = (_zz_when_BankedScratchMemory_l242_15 == 3'b110);
  assign when_BankedScratchMemory_l242_127 = (_zz_when_BankedScratchMemory_l242_15 == 3'b111);
  assign _zz_when_BankedScratchMemory_l242_16 = io_writeAddr_16[2 : 0];
  assign _zz_io_write_addr_16 = io_writeAddr_16[10 : 3];
  assign when_BankedScratchMemory_l242_128 = (_zz_when_BankedScratchMemory_l242_16 == 3'b000);
  assign when_BankedScratchMemory_l242_129 = (_zz_when_BankedScratchMemory_l242_16 == 3'b001);
  assign when_BankedScratchMemory_l242_130 = (_zz_when_BankedScratchMemory_l242_16 == 3'b010);
  assign when_BankedScratchMemory_l242_131 = (_zz_when_BankedScratchMemory_l242_16 == 3'b011);
  assign when_BankedScratchMemory_l242_132 = (_zz_when_BankedScratchMemory_l242_16 == 3'b100);
  assign when_BankedScratchMemory_l242_133 = (_zz_when_BankedScratchMemory_l242_16 == 3'b101);
  assign when_BankedScratchMemory_l242_134 = (_zz_when_BankedScratchMemory_l242_16 == 3'b110);
  assign when_BankedScratchMemory_l242_135 = (_zz_when_BankedScratchMemory_l242_16 == 3'b111);
  assign _zz_when_BankedScratchMemory_l242_17 = io_writeAddr_17[2 : 0];
  assign _zz_io_write_addr_17 = io_writeAddr_17[10 : 3];
  assign when_BankedScratchMemory_l242_136 = (_zz_when_BankedScratchMemory_l242_17 == 3'b000);
  assign when_BankedScratchMemory_l242_137 = (_zz_when_BankedScratchMemory_l242_17 == 3'b001);
  assign when_BankedScratchMemory_l242_138 = (_zz_when_BankedScratchMemory_l242_17 == 3'b010);
  assign when_BankedScratchMemory_l242_139 = (_zz_when_BankedScratchMemory_l242_17 == 3'b011);
  assign when_BankedScratchMemory_l242_140 = (_zz_when_BankedScratchMemory_l242_17 == 3'b100);
  assign when_BankedScratchMemory_l242_141 = (_zz_when_BankedScratchMemory_l242_17 == 3'b101);
  assign when_BankedScratchMemory_l242_142 = (_zz_when_BankedScratchMemory_l242_17 == 3'b110);
  assign when_BankedScratchMemory_l242_143 = (_zz_when_BankedScratchMemory_l242_17 == 3'b111);
  assign _zz_when_BankedScratchMemory_l242_18 = io_writeAddr_18[2 : 0];
  assign _zz_io_write_addr_18 = io_writeAddr_18[10 : 3];
  assign when_BankedScratchMemory_l242_144 = (_zz_when_BankedScratchMemory_l242_18 == 3'b000);
  assign when_BankedScratchMemory_l242_145 = (_zz_when_BankedScratchMemory_l242_18 == 3'b001);
  assign when_BankedScratchMemory_l242_146 = (_zz_when_BankedScratchMemory_l242_18 == 3'b010);
  assign when_BankedScratchMemory_l242_147 = (_zz_when_BankedScratchMemory_l242_18 == 3'b011);
  assign when_BankedScratchMemory_l242_148 = (_zz_when_BankedScratchMemory_l242_18 == 3'b100);
  assign when_BankedScratchMemory_l242_149 = (_zz_when_BankedScratchMemory_l242_18 == 3'b101);
  assign when_BankedScratchMemory_l242_150 = (_zz_when_BankedScratchMemory_l242_18 == 3'b110);
  assign when_BankedScratchMemory_l242_151 = (_zz_when_BankedScratchMemory_l242_18 == 3'b111);
  assign _zz_when_BankedScratchMemory_l242_19 = io_writeAddr_19[2 : 0];
  assign _zz_io_write_addr_19 = io_writeAddr_19[10 : 3];
  assign when_BankedScratchMemory_l242_152 = (_zz_when_BankedScratchMemory_l242_19 == 3'b000);
  assign when_BankedScratchMemory_l242_153 = (_zz_when_BankedScratchMemory_l242_19 == 3'b001);
  assign when_BankedScratchMemory_l242_154 = (_zz_when_BankedScratchMemory_l242_19 == 3'b010);
  assign when_BankedScratchMemory_l242_155 = (_zz_when_BankedScratchMemory_l242_19 == 3'b011);
  assign when_BankedScratchMemory_l242_156 = (_zz_when_BankedScratchMemory_l242_19 == 3'b100);
  assign when_BankedScratchMemory_l242_157 = (_zz_when_BankedScratchMemory_l242_19 == 3'b101);
  assign when_BankedScratchMemory_l242_158 = (_zz_when_BankedScratchMemory_l242_19 == 3'b110);
  assign when_BankedScratchMemory_l242_159 = (_zz_when_BankedScratchMemory_l242_19 == 3'b111);
  assign _zz_when_BankedScratchMemory_l242_20 = io_writeAddr_20[2 : 0];
  assign _zz_io_write_addr_20 = io_writeAddr_20[10 : 3];
  assign when_BankedScratchMemory_l242_160 = (_zz_when_BankedScratchMemory_l242_20 == 3'b000);
  assign when_BankedScratchMemory_l242_161 = (_zz_when_BankedScratchMemory_l242_20 == 3'b001);
  assign when_BankedScratchMemory_l242_162 = (_zz_when_BankedScratchMemory_l242_20 == 3'b010);
  assign when_BankedScratchMemory_l242_163 = (_zz_when_BankedScratchMemory_l242_20 == 3'b011);
  assign when_BankedScratchMemory_l242_164 = (_zz_when_BankedScratchMemory_l242_20 == 3'b100);
  assign when_BankedScratchMemory_l242_165 = (_zz_when_BankedScratchMemory_l242_20 == 3'b101);
  assign when_BankedScratchMemory_l242_166 = (_zz_when_BankedScratchMemory_l242_20 == 3'b110);
  assign when_BankedScratchMemory_l242_167 = (_zz_when_BankedScratchMemory_l242_20 == 3'b111);
  assign _zz_when_BankedScratchMemory_l242_21 = io_writeAddr_21[2 : 0];
  assign _zz_io_write_addr_21 = io_writeAddr_21[10 : 3];
  assign when_BankedScratchMemory_l242_168 = (_zz_when_BankedScratchMemory_l242_21 == 3'b000);
  assign when_BankedScratchMemory_l242_169 = (_zz_when_BankedScratchMemory_l242_21 == 3'b001);
  assign when_BankedScratchMemory_l242_170 = (_zz_when_BankedScratchMemory_l242_21 == 3'b010);
  assign when_BankedScratchMemory_l242_171 = (_zz_when_BankedScratchMemory_l242_21 == 3'b011);
  assign when_BankedScratchMemory_l242_172 = (_zz_when_BankedScratchMemory_l242_21 == 3'b100);
  assign when_BankedScratchMemory_l242_173 = (_zz_when_BankedScratchMemory_l242_21 == 3'b101);
  assign when_BankedScratchMemory_l242_174 = (_zz_when_BankedScratchMemory_l242_21 == 3'b110);
  assign when_BankedScratchMemory_l242_175 = (_zz_when_BankedScratchMemory_l242_21 == 3'b111);
  assign _zz_when_BankedScratchMemory_l242_22 = io_writeAddr_22[2 : 0];
  assign _zz_io_write_addr_22 = io_writeAddr_22[10 : 3];
  assign when_BankedScratchMemory_l242_176 = (_zz_when_BankedScratchMemory_l242_22 == 3'b000);
  assign when_BankedScratchMemory_l242_177 = (_zz_when_BankedScratchMemory_l242_22 == 3'b001);
  assign when_BankedScratchMemory_l242_178 = (_zz_when_BankedScratchMemory_l242_22 == 3'b010);
  assign when_BankedScratchMemory_l242_179 = (_zz_when_BankedScratchMemory_l242_22 == 3'b011);
  assign when_BankedScratchMemory_l242_180 = (_zz_when_BankedScratchMemory_l242_22 == 3'b100);
  assign when_BankedScratchMemory_l242_181 = (_zz_when_BankedScratchMemory_l242_22 == 3'b101);
  assign when_BankedScratchMemory_l242_182 = (_zz_when_BankedScratchMemory_l242_22 == 3'b110);
  assign when_BankedScratchMemory_l242_183 = (_zz_when_BankedScratchMemory_l242_22 == 3'b111);
  assign _zz_when_BankedScratchMemory_l242_23 = io_writeAddr_23[2 : 0];
  assign _zz_io_write_addr_23 = io_writeAddr_23[10 : 3];
  assign when_BankedScratchMemory_l242_184 = (_zz_when_BankedScratchMemory_l242_23 == 3'b000);
  assign when_BankedScratchMemory_l242_185 = (_zz_when_BankedScratchMemory_l242_23 == 3'b001);
  assign when_BankedScratchMemory_l242_186 = (_zz_when_BankedScratchMemory_l242_23 == 3'b010);
  assign when_BankedScratchMemory_l242_187 = (_zz_when_BankedScratchMemory_l242_23 == 3'b011);
  assign when_BankedScratchMemory_l242_188 = (_zz_when_BankedScratchMemory_l242_23 == 3'b100);
  assign when_BankedScratchMemory_l242_189 = (_zz_when_BankedScratchMemory_l242_23 == 3'b101);
  assign when_BankedScratchMemory_l242_190 = (_zz_when_BankedScratchMemory_l242_23 == 3'b110);
  assign when_BankedScratchMemory_l242_191 = (_zz_when_BankedScratchMemory_l242_23 == 3'b111);
  assign _zz_when_BankedScratchMemory_l242_24 = io_writeAddr_24[2 : 0];
  assign _zz_io_write_addr_24 = io_writeAddr_24[10 : 3];
  assign when_BankedScratchMemory_l242_192 = (_zz_when_BankedScratchMemory_l242_24 == 3'b000);
  assign when_BankedScratchMemory_l242_193 = (_zz_when_BankedScratchMemory_l242_24 == 3'b001);
  assign when_BankedScratchMemory_l242_194 = (_zz_when_BankedScratchMemory_l242_24 == 3'b010);
  assign when_BankedScratchMemory_l242_195 = (_zz_when_BankedScratchMemory_l242_24 == 3'b011);
  assign when_BankedScratchMemory_l242_196 = (_zz_when_BankedScratchMemory_l242_24 == 3'b100);
  assign when_BankedScratchMemory_l242_197 = (_zz_when_BankedScratchMemory_l242_24 == 3'b101);
  assign when_BankedScratchMemory_l242_198 = (_zz_when_BankedScratchMemory_l242_24 == 3'b110);
  assign when_BankedScratchMemory_l242_199 = (_zz_when_BankedScratchMemory_l242_24 == 3'b111);
  assign _zz_when_BankedScratchMemory_l242_25 = io_writeAddr_25[2 : 0];
  assign _zz_io_write_addr_25 = io_writeAddr_25[10 : 3];
  assign when_BankedScratchMemory_l242_200 = (_zz_when_BankedScratchMemory_l242_25 == 3'b000);
  assign when_BankedScratchMemory_l242_201 = (_zz_when_BankedScratchMemory_l242_25 == 3'b001);
  assign when_BankedScratchMemory_l242_202 = (_zz_when_BankedScratchMemory_l242_25 == 3'b010);
  assign when_BankedScratchMemory_l242_203 = (_zz_when_BankedScratchMemory_l242_25 == 3'b011);
  assign when_BankedScratchMemory_l242_204 = (_zz_when_BankedScratchMemory_l242_25 == 3'b100);
  assign when_BankedScratchMemory_l242_205 = (_zz_when_BankedScratchMemory_l242_25 == 3'b101);
  assign when_BankedScratchMemory_l242_206 = (_zz_when_BankedScratchMemory_l242_25 == 3'b110);
  assign when_BankedScratchMemory_l242_207 = (_zz_when_BankedScratchMemory_l242_25 == 3'b111);
  assign _zz_when_BankedScratchMemory_l242_26 = io_writeAddr_26[2 : 0];
  assign _zz_io_write_addr_26 = io_writeAddr_26[10 : 3];
  assign when_BankedScratchMemory_l242_208 = (_zz_when_BankedScratchMemory_l242_26 == 3'b000);
  assign when_BankedScratchMemory_l242_209 = (_zz_when_BankedScratchMemory_l242_26 == 3'b001);
  assign when_BankedScratchMemory_l242_210 = (_zz_when_BankedScratchMemory_l242_26 == 3'b010);
  assign when_BankedScratchMemory_l242_211 = (_zz_when_BankedScratchMemory_l242_26 == 3'b011);
  assign when_BankedScratchMemory_l242_212 = (_zz_when_BankedScratchMemory_l242_26 == 3'b100);
  assign when_BankedScratchMemory_l242_213 = (_zz_when_BankedScratchMemory_l242_26 == 3'b101);
  assign when_BankedScratchMemory_l242_214 = (_zz_when_BankedScratchMemory_l242_26 == 3'b110);
  assign when_BankedScratchMemory_l242_215 = (_zz_when_BankedScratchMemory_l242_26 == 3'b111);
  assign _zz_when_BankedScratchMemory_l242_27 = io_writeAddr_27[2 : 0];
  assign _zz_io_write_addr_27 = io_writeAddr_27[10 : 3];
  assign when_BankedScratchMemory_l242_216 = (_zz_when_BankedScratchMemory_l242_27 == 3'b000);
  assign when_BankedScratchMemory_l242_217 = (_zz_when_BankedScratchMemory_l242_27 == 3'b001);
  assign when_BankedScratchMemory_l242_218 = (_zz_when_BankedScratchMemory_l242_27 == 3'b010);
  assign when_BankedScratchMemory_l242_219 = (_zz_when_BankedScratchMemory_l242_27 == 3'b011);
  assign when_BankedScratchMemory_l242_220 = (_zz_when_BankedScratchMemory_l242_27 == 3'b100);
  assign when_BankedScratchMemory_l242_221 = (_zz_when_BankedScratchMemory_l242_27 == 3'b101);
  assign when_BankedScratchMemory_l242_222 = (_zz_when_BankedScratchMemory_l242_27 == 3'b110);
  assign when_BankedScratchMemory_l242_223 = (_zz_when_BankedScratchMemory_l242_27 == 3'b111);

endmodule

module DecodeUnit (
  input  wire [255:0]  io_bundle,
  input  wire          io_valid,
  output wire          io_aluSlots_0_valid,
  output wire [3:0]    io_aluSlots_0_opcode,
  output wire [10:0]   io_aluSlots_0_dest,
  output wire [10:0]   io_aluSlots_0_src1,
  output wire [10:0]   io_aluSlots_0_src2,
  output wire          io_valuSlots_0_valid,
  output wire [3:0]    io_valuSlots_0_opcode,
  output wire [10:0]   io_valuSlots_0_destBase,
  output wire [10:0]   io_valuSlots_0_src1Base,
  output wire [10:0]   io_valuSlots_0_src2Base,
  output wire [10:0]   io_valuSlots_0_src3Base,
  output wire          io_loadSlots_0_valid,
  output wire [2:0]    io_loadSlots_0_opcode,
  output wire [10:0]   io_loadSlots_0_dest,
  output wire [10:0]   io_loadSlots_0_addrReg,
  output wire [2:0]    io_loadSlots_0_offset,
  output wire [31:0]   io_loadSlots_0_immediate,
  output wire          io_storeSlots_0_valid,
  output wire [1:0]    io_storeSlots_0_opcode,
  output wire [10:0]   io_storeSlots_0_addrReg,
  output wire [10:0]   io_storeSlots_0_srcReg,
  output wire          io_flowSlot_valid,
  output wire [3:0]    io_flowSlot_opcode,
  output wire [10:0]   io_flowSlot_dest,
  output wire [10:0]   io_flowSlot_operandA,
  output wire [10:0]   io_flowSlot_operandB,
  output wire [9:0]    io_flowSlot_immediate
);

  wire       [39:0]   _zz_io_aluSlots_0_valid;
  wire       [55:0]   _zz_io_valuSlots_0_valid;
  wire       [47:0]   _zz_io_loadSlots_0_valid;
  wire       [27:0]   _zz_io_storeSlots_0_valid;
  wire       [47:0]   _zz_io_flowSlot_valid;

  assign _zz_io_aluSlots_0_valid = io_bundle[39 : 0];
  assign io_aluSlots_0_valid = (_zz_io_aluSlots_0_valid[39] && io_valid);
  assign io_aluSlots_0_opcode = _zz_io_aluSlots_0_valid[38 : 35];
  assign io_aluSlots_0_dest = _zz_io_aluSlots_0_valid[34 : 24];
  assign io_aluSlots_0_src1 = _zz_io_aluSlots_0_valid[23 : 13];
  assign io_aluSlots_0_src2 = _zz_io_aluSlots_0_valid[12 : 2];
  assign _zz_io_valuSlots_0_valid = io_bundle[95 : 40];
  assign io_valuSlots_0_valid = (_zz_io_valuSlots_0_valid[55] && io_valid);
  assign io_valuSlots_0_opcode = _zz_io_valuSlots_0_valid[54 : 51];
  assign io_valuSlots_0_destBase = _zz_io_valuSlots_0_valid[50 : 40];
  assign io_valuSlots_0_src1Base = _zz_io_valuSlots_0_valid[39 : 29];
  assign io_valuSlots_0_src2Base = _zz_io_valuSlots_0_valid[28 : 18];
  assign io_valuSlots_0_src3Base = _zz_io_valuSlots_0_valid[17 : 7];
  assign _zz_io_loadSlots_0_valid = io_bundle[143 : 96];
  assign io_loadSlots_0_valid = (_zz_io_loadSlots_0_valid[47] && io_valid);
  assign io_loadSlots_0_opcode = _zz_io_loadSlots_0_valid[46 : 44];
  assign io_loadSlots_0_dest = _zz_io_loadSlots_0_valid[43 : 33];
  assign io_loadSlots_0_addrReg = _zz_io_loadSlots_0_valid[32 : 22];
  assign io_loadSlots_0_offset = _zz_io_loadSlots_0_valid[21 : 19];
  assign io_loadSlots_0_immediate = _zz_io_loadSlots_0_valid[31 : 0];
  assign _zz_io_storeSlots_0_valid = io_bundle[171 : 144];
  assign io_storeSlots_0_valid = (_zz_io_storeSlots_0_valid[27] && io_valid);
  assign io_storeSlots_0_opcode = _zz_io_storeSlots_0_valid[26 : 25];
  assign io_storeSlots_0_addrReg = _zz_io_storeSlots_0_valid[24 : 14];
  assign io_storeSlots_0_srcReg = _zz_io_storeSlots_0_valid[13 : 3];
  assign _zz_io_flowSlot_valid = io_bundle[219 : 172];
  assign io_flowSlot_valid = (_zz_io_flowSlot_valid[47] && io_valid);
  assign io_flowSlot_opcode = _zz_io_flowSlot_valid[46 : 43];
  assign io_flowSlot_dest = _zz_io_flowSlot_valid[42 : 32];
  assign io_flowSlot_operandA = _zz_io_flowSlot_valid[31 : 21];
  assign io_flowSlot_operandB = _zz_io_flowSlot_valid[20 : 10];
  assign io_flowSlot_immediate = _zz_io_flowSlot_valid[9 : 0];

endmodule

module FetchUnit (
  output wire [9:0]    io_imemAddr,
  input  wire [255:0]  io_imemData,
  output wire [255:0]  io_exBundle,
  output wire          io_exValid,
  input  wire          io_jump_valid,
  input  wire [9:0]    io_jump_payload,
  input  wire          io_halt,
  input  wire          io_start,
  input  wire          io_stall,
  output wire [9:0]    io_pc,
  output wire          io_running,
  output wire          io_halted,
  input  wire          clk,
  input  wire          reset
);
  localparam CoreState_IDLE = 2'd0;
  localparam CoreState_RUNNING = 2'd1;
  localparam CoreState_HALTED = 2'd2;

  reg        [1:0]    state;
  reg        [9:0]    pc;
  wire                cycleActive;
  reg        [255:0]  exBundleReg;
  reg                 exValidReg;
  wire                when_FetchUnit_l80;
  `ifndef SYNTHESIS
  reg [55:0] state_string;
  `endif


  `ifndef SYNTHESIS
  always @(*) begin
    case(state)
      CoreState_IDLE : state_string = "IDLE   ";
      CoreState_RUNNING : state_string = "RUNNING";
      CoreState_HALTED : state_string = "HALTED ";
      default : state_string = "???????";
    endcase
  end
  `endif

  assign cycleActive = (state == CoreState_RUNNING);
  assign io_imemAddr = pc;
  assign when_FetchUnit_l80 = (! io_stall);
  assign io_exBundle = exBundleReg;
  assign io_exValid = exValidReg;
  assign io_pc = pc;
  assign io_running = cycleActive;
  assign io_halted = (state == CoreState_HALTED);
  always @(posedge clk) begin
    if(reset) begin
      state <= CoreState_IDLE;
      pc <= 10'h0;
      exBundleReg <= 256'h0;
      exValidReg <= 1'b0;
    end else begin
      case(state)
        CoreState_IDLE : begin
          if(io_start) begin
            state <= CoreState_RUNNING;
            pc <= 10'h0;
          end
        end
        CoreState_RUNNING : begin
          if(io_halt) begin
            state <= CoreState_HALTED;
          end
        end
        default : begin
          if(io_start) begin
            state <= CoreState_RUNNING;
            pc <= 10'h0;
          end
        end
      endcase
      if(when_FetchUnit_l80) begin
        if(cycleActive) begin
          if(io_jump_valid) begin
            pc <= io_jump_payload;
            exValidReg <= 1'b0;
            exBundleReg <= 256'h0;
          end else begin
            if(io_halt) begin
              exValidReg <= 1'b0;
            end else begin
              exBundleReg <= io_imemData;
              exValidReg <= 1'b1;
              pc <= (pc + 10'h001);
            end
          end
        end else begin
          exValidReg <= 1'b0;
        end
      end
    end
  end


endmodule

module InstructionMemory (
  input  wire [9:0]    io_fetchAddr,
  output wire [255:0]  io_fetchData,
  input  wire          io_write_valid,
  input  wire [9:0]    io_write_payload_addr,
  input  wire [255:0]  io_write_payload_data,
  input  wire          clk,
  input  wire          reset
);

  reg        [255:0]  mem_spinal_port0;
  wire                _zz_mem_port;
  wire                _zz_io_fetchData;
  reg                 _zz_1;
  reg [255:0] mem [0:1023];

  assign _zz_io_fetchData = 1'b1;
  always @(posedge clk) begin
    if(_zz_io_fetchData) begin
      mem_spinal_port0 <= mem[io_fetchAddr];
    end
  end

  always @(posedge clk) begin
    if(_zz_1) begin
      mem[io_write_payload_addr] <= io_write_payload_data;
    end
  end

  always @(*) begin
    _zz_1 = 1'b0;
    if(io_write_valid) begin
      _zz_1 = 1'b1;
    end
  end

  assign io_fetchData = mem_spinal_port0;

endmodule

module StreamFifoLowLatency (
  input  wire          io_push_valid,
  output wire          io_push_ready,
  input  wire [0:0]    io_push_payload,
  output wire          io_pop_valid,
  input  wire          io_pop_ready,
  output wire [0:0]    io_pop_payload,
  input  wire          io_flush,
  output wire [2:0]    io_occupancy,
  output wire [2:0]    io_availability,
  input  wire          clk,
  input  wire          reset
);

  wire                fifo_io_push_ready;
  wire                fifo_io_pop_valid;
  wire       [0:0]    fifo_io_pop_payload;
  wire       [2:0]    fifo_io_occupancy;
  wire       [2:0]    fifo_io_availability;

  StreamFifo fifo (
    .io_push_valid   (io_push_valid            ), //i
    .io_push_ready   (fifo_io_push_ready       ), //o
    .io_push_payload (io_push_payload          ), //i
    .io_pop_valid    (fifo_io_pop_valid        ), //o
    .io_pop_ready    (io_pop_ready             ), //i
    .io_pop_payload  (fifo_io_pop_payload      ), //o
    .io_flush        (io_flush                 ), //i
    .io_occupancy    (fifo_io_occupancy[2:0]   ), //o
    .io_availability (fifo_io_availability[2:0]), //o
    .clk             (clk                      ), //i
    .reset           (reset                    )  //i
  );
  assign io_push_ready = fifo_io_push_ready;
  assign io_pop_valid = fifo_io_pop_valid;
  assign io_pop_payload = fifo_io_pop_payload;
  assign io_occupancy = fifo_io_occupancy;
  assign io_availability = fifo_io_availability;

endmodule

module StreamArbiter (
  input  wire          io_inputs_0_valid,
  output wire          io_inputs_0_ready,
  input  wire [15:0]   io_inputs_0_payload_addr,
  input  wire [4:0]    io_inputs_0_payload_id,
  input  wire [7:0]    io_inputs_0_payload_len,
  input  wire [2:0]    io_inputs_0_payload_size,
  input  wire [1:0]    io_inputs_0_payload_burst,
  input  wire          io_inputs_0_payload_write,
  input  wire          io_inputs_1_valid,
  output wire          io_inputs_1_ready,
  input  wire [15:0]   io_inputs_1_payload_addr,
  input  wire [4:0]    io_inputs_1_payload_id,
  input  wire [7:0]    io_inputs_1_payload_len,
  input  wire [2:0]    io_inputs_1_payload_size,
  input  wire [1:0]    io_inputs_1_payload_burst,
  input  wire          io_inputs_1_payload_write,
  input  wire          io_inputs_2_valid,
  output wire          io_inputs_2_ready,
  input  wire [15:0]   io_inputs_2_payload_addr,
  input  wire [4:0]    io_inputs_2_payload_id,
  input  wire [7:0]    io_inputs_2_payload_len,
  input  wire [2:0]    io_inputs_2_payload_size,
  input  wire [1:0]    io_inputs_2_payload_burst,
  input  wire          io_inputs_2_payload_write,
  input  wire          io_inputs_3_valid,
  output wire          io_inputs_3_ready,
  input  wire [15:0]   io_inputs_3_payload_addr,
  input  wire [4:0]    io_inputs_3_payload_id,
  input  wire [7:0]    io_inputs_3_payload_len,
  input  wire [2:0]    io_inputs_3_payload_size,
  input  wire [1:0]    io_inputs_3_payload_burst,
  input  wire          io_inputs_3_payload_write,
  output wire          io_output_valid,
  input  wire          io_output_ready,
  output wire [15:0]   io_output_payload_addr,
  output wire [4:0]    io_output_payload_id,
  output wire [7:0]    io_output_payload_len,
  output wire [2:0]    io_output_payload_size,
  output wire [1:0]    io_output_payload_burst,
  output wire          io_output_payload_write,
  output wire [1:0]    io_chosen,
  output wire [3:0]    io_chosenOH,
  input  wire          clk,
  input  wire          reset
);

  wire       [7:0]    _zz__zz_maskProposal_0_2;
  wire       [7:0]    _zz__zz_maskProposal_0_2_1;
  wire       [3:0]    _zz__zz_maskProposal_0_2_2;
  reg        [15:0]   _zz_io_output_payload_addr_3;
  reg        [4:0]    _zz_io_output_payload_id;
  reg        [7:0]    _zz_io_output_payload_len;
  reg        [2:0]    _zz_io_output_payload_size;
  reg        [1:0]    _zz_io_output_payload_burst;
  reg                 _zz_io_output_payload_write;
  reg                 locked;
  wire                maskProposal_0;
  wire                maskProposal_1;
  wire                maskProposal_2;
  wire                maskProposal_3;
  reg                 maskLocked_0;
  reg                 maskLocked_1;
  reg                 maskLocked_2;
  reg                 maskLocked_3;
  wire                maskRouted_0;
  wire                maskRouted_1;
  wire                maskRouted_2;
  wire                maskRouted_3;
  wire       [3:0]    _zz_maskProposal_0;
  wire       [7:0]    _zz_maskProposal_0_1;
  wire       [7:0]    _zz_maskProposal_0_2;
  wire       [3:0]    _zz_maskProposal_0_3;
  wire                io_output_fire;
  wire                _zz_io_output_payload_addr;
  wire                _zz_io_output_payload_addr_1;
  wire       [1:0]    _zz_io_output_payload_addr_2;
  wire                _zz_io_chosen;
  wire                _zz_io_chosen_1;
  wire                _zz_io_chosen_2;

  assign _zz__zz_maskProposal_0_2 = (_zz_maskProposal_0_1 - _zz__zz_maskProposal_0_2_1);
  assign _zz__zz_maskProposal_0_2_2 = {maskLocked_2,{maskLocked_1,{maskLocked_0,maskLocked_3}}};
  assign _zz__zz_maskProposal_0_2_1 = {4'd0, _zz__zz_maskProposal_0_2_2};
  always @(*) begin
    case(_zz_io_output_payload_addr_2)
      2'b00 : begin
        _zz_io_output_payload_addr_3 = io_inputs_0_payload_addr;
        _zz_io_output_payload_id = io_inputs_0_payload_id;
        _zz_io_output_payload_len = io_inputs_0_payload_len;
        _zz_io_output_payload_size = io_inputs_0_payload_size;
        _zz_io_output_payload_burst = io_inputs_0_payload_burst;
        _zz_io_output_payload_write = io_inputs_0_payload_write;
      end
      2'b01 : begin
        _zz_io_output_payload_addr_3 = io_inputs_1_payload_addr;
        _zz_io_output_payload_id = io_inputs_1_payload_id;
        _zz_io_output_payload_len = io_inputs_1_payload_len;
        _zz_io_output_payload_size = io_inputs_1_payload_size;
        _zz_io_output_payload_burst = io_inputs_1_payload_burst;
        _zz_io_output_payload_write = io_inputs_1_payload_write;
      end
      2'b10 : begin
        _zz_io_output_payload_addr_3 = io_inputs_2_payload_addr;
        _zz_io_output_payload_id = io_inputs_2_payload_id;
        _zz_io_output_payload_len = io_inputs_2_payload_len;
        _zz_io_output_payload_size = io_inputs_2_payload_size;
        _zz_io_output_payload_burst = io_inputs_2_payload_burst;
        _zz_io_output_payload_write = io_inputs_2_payload_write;
      end
      default : begin
        _zz_io_output_payload_addr_3 = io_inputs_3_payload_addr;
        _zz_io_output_payload_id = io_inputs_3_payload_id;
        _zz_io_output_payload_len = io_inputs_3_payload_len;
        _zz_io_output_payload_size = io_inputs_3_payload_size;
        _zz_io_output_payload_burst = io_inputs_3_payload_burst;
        _zz_io_output_payload_write = io_inputs_3_payload_write;
      end
    endcase
  end

  assign maskRouted_0 = (locked ? maskLocked_0 : maskProposal_0);
  assign maskRouted_1 = (locked ? maskLocked_1 : maskProposal_1);
  assign maskRouted_2 = (locked ? maskLocked_2 : maskProposal_2);
  assign maskRouted_3 = (locked ? maskLocked_3 : maskProposal_3);
  assign _zz_maskProposal_0 = {io_inputs_3_valid,{io_inputs_2_valid,{io_inputs_1_valid,io_inputs_0_valid}}};
  assign _zz_maskProposal_0_1 = {_zz_maskProposal_0,_zz_maskProposal_0};
  assign _zz_maskProposal_0_2 = (_zz_maskProposal_0_1 & (~ _zz__zz_maskProposal_0_2));
  assign _zz_maskProposal_0_3 = (_zz_maskProposal_0_2[7 : 4] | _zz_maskProposal_0_2[3 : 0]);
  assign maskProposal_0 = _zz_maskProposal_0_3[0];
  assign maskProposal_1 = _zz_maskProposal_0_3[1];
  assign maskProposal_2 = _zz_maskProposal_0_3[2];
  assign maskProposal_3 = _zz_maskProposal_0_3[3];
  assign io_output_fire = (io_output_valid && io_output_ready);
  assign io_output_valid = ((((io_inputs_0_valid && maskRouted_0) || (io_inputs_1_valid && maskRouted_1)) || (io_inputs_2_valid && maskRouted_2)) || (io_inputs_3_valid && maskRouted_3));
  assign _zz_io_output_payload_addr = (maskRouted_1 || maskRouted_3);
  assign _zz_io_output_payload_addr_1 = (maskRouted_2 || maskRouted_3);
  assign _zz_io_output_payload_addr_2 = {_zz_io_output_payload_addr_1,_zz_io_output_payload_addr};
  assign io_output_payload_addr = _zz_io_output_payload_addr_3;
  assign io_output_payload_id = _zz_io_output_payload_id;
  assign io_output_payload_len = _zz_io_output_payload_len;
  assign io_output_payload_size = _zz_io_output_payload_size;
  assign io_output_payload_burst = _zz_io_output_payload_burst;
  assign io_output_payload_write = _zz_io_output_payload_write;
  assign io_inputs_0_ready = (maskRouted_0 && io_output_ready);
  assign io_inputs_1_ready = (maskRouted_1 && io_output_ready);
  assign io_inputs_2_ready = (maskRouted_2 && io_output_ready);
  assign io_inputs_3_ready = (maskRouted_3 && io_output_ready);
  assign io_chosenOH = {maskRouted_3,{maskRouted_2,{maskRouted_1,maskRouted_0}}};
  assign _zz_io_chosen = io_chosenOH[3];
  assign _zz_io_chosen_1 = (io_chosenOH[1] || _zz_io_chosen);
  assign _zz_io_chosen_2 = (io_chosenOH[2] || _zz_io_chosen);
  assign io_chosen = {_zz_io_chosen_2,_zz_io_chosen_1};
  always @(posedge clk) begin
    if(reset) begin
      locked <= 1'b0;
      maskLocked_0 <= 1'b0;
      maskLocked_1 <= 1'b0;
      maskLocked_2 <= 1'b0;
      maskLocked_3 <= 1'b1;
    end else begin
      if(io_output_valid) begin
        maskLocked_0 <= maskRouted_0;
        maskLocked_1 <= maskRouted_1;
        maskLocked_2 <= maskRouted_2;
        maskLocked_3 <= maskRouted_3;
      end
      if(io_output_valid) begin
        locked <= 1'b1;
      end
      if(io_output_fire) begin
        locked <= 1'b0;
      end
    end
  end


endmodule

//Axi4WriteOnlyErrorSlave replaced by Axi4WriteOnlyErrorSlave_1

//Axi4ReadOnlyErrorSlave replaced by Axi4ReadOnlyErrorSlave_1

module Axi4WriteOnlyErrorSlave_1 (
  input  wire          io_axi_aw_valid,
  output wire          io_axi_aw_ready,
  input  wire [31:0]   io_axi_aw_payload_addr,
  input  wire [3:0]    io_axi_aw_payload_id,
  input  wire [7:0]    io_axi_aw_payload_len,
  input  wire [2:0]    io_axi_aw_payload_size,
  input  wire [1:0]    io_axi_aw_payload_burst,
  input  wire          io_axi_w_valid,
  output wire          io_axi_w_ready,
  input  wire [31:0]   io_axi_w_payload_data,
  input  wire [3:0]    io_axi_w_payload_strb,
  input  wire          io_axi_w_payload_last,
  output wire          io_axi_b_valid,
  input  wire          io_axi_b_ready,
  output wire [3:0]    io_axi_b_payload_id,
  output wire [1:0]    io_axi_b_payload_resp,
  input  wire          clk,
  input  wire          reset
);

  reg                 consumeData;
  reg                 sendRsp;
  reg        [3:0]    id;
  wire                io_axi_aw_fire;
  wire                io_axi_w_fire;
  wire                when_Axi4ErrorSlave_l24;
  wire                io_axi_b_fire;

  assign io_axi_aw_ready = (! (consumeData || sendRsp));
  assign io_axi_aw_fire = (io_axi_aw_valid && io_axi_aw_ready);
  assign io_axi_w_ready = consumeData;
  assign io_axi_w_fire = (io_axi_w_valid && io_axi_w_ready);
  assign when_Axi4ErrorSlave_l24 = (io_axi_w_fire && io_axi_w_payload_last);
  assign io_axi_b_valid = sendRsp;
  assign io_axi_b_payload_resp = 2'b11;
  assign io_axi_b_payload_id = id;
  assign io_axi_b_fire = (io_axi_b_valid && io_axi_b_ready);
  always @(posedge clk) begin
    if(reset) begin
      consumeData <= 1'b0;
      sendRsp <= 1'b0;
    end else begin
      if(io_axi_aw_fire) begin
        consumeData <= 1'b1;
      end
      if(when_Axi4ErrorSlave_l24) begin
        consumeData <= 1'b0;
        sendRsp <= 1'b1;
      end
      if(io_axi_b_fire) begin
        sendRsp <= 1'b0;
      end
    end
  end

  always @(posedge clk) begin
    if(io_axi_aw_fire) begin
      id <= io_axi_aw_payload_id;
    end
  end


endmodule

module Axi4ReadOnlyErrorSlave_1 (
  input  wire          io_axi_ar_valid,
  output wire          io_axi_ar_ready,
  input  wire [31:0]   io_axi_ar_payload_addr,
  input  wire [3:0]    io_axi_ar_payload_id,
  input  wire [7:0]    io_axi_ar_payload_len,
  input  wire [2:0]    io_axi_ar_payload_size,
  input  wire [1:0]    io_axi_ar_payload_burst,
  output wire          io_axi_r_valid,
  input  wire          io_axi_r_ready,
  output wire [31:0]   io_axi_r_payload_data,
  output wire [3:0]    io_axi_r_payload_id,
  output wire [1:0]    io_axi_r_payload_resp,
  output wire          io_axi_r_payload_last,
  input  wire          clk,
  input  wire          reset
);

  reg                 sendRsp;
  reg        [3:0]    id;
  reg        [7:0]    remaining;
  wire                remainingZero;
  wire                io_axi_ar_fire;

  assign remainingZero = (remaining == 8'h0);
  assign io_axi_ar_ready = (! sendRsp);
  assign io_axi_ar_fire = (io_axi_ar_valid && io_axi_ar_ready);
  assign io_axi_r_valid = sendRsp;
  assign io_axi_r_payload_id = id;
  assign io_axi_r_payload_resp = 2'b11;
  assign io_axi_r_payload_last = remainingZero;
  always @(posedge clk) begin
    if(reset) begin
      sendRsp <= 1'b0;
    end else begin
      if(io_axi_ar_fire) begin
        sendRsp <= 1'b1;
      end
      if(sendRsp) begin
        if(io_axi_r_ready) begin
          if(remainingZero) begin
            sendRsp <= 1'b0;
          end
        end
      end
    end
  end

  always @(posedge clk) begin
    if(io_axi_ar_fire) begin
      remaining <= io_axi_ar_payload_len;
      id <= io_axi_ar_payload_id;
    end
    if(sendRsp) begin
      if(io_axi_r_ready) begin
        remaining <= (remaining - 8'h01);
      end
    end
  end


endmodule

//UnsignedDivider_7 replaced by UnsignedDivider_8

//UnsignedDivider_6 replaced by UnsignedDivider_8

//UnsignedDivider_5 replaced by UnsignedDivider_8

//UnsignedDivider_4 replaced by UnsignedDivider_8

//UnsignedDivider_3 replaced by UnsignedDivider_8

//UnsignedDivider_2 replaced by UnsignedDivider_8

//UnsignedDivider_1 replaced by UnsignedDivider_8

//UnsignedDivider replaced by UnsignedDivider_8

module UnsignedDivider_8 (
  input  wire          io_start,
  input  wire [31:0]   io_dividend,
  input  wire [31:0]   io_divisor,
  output wire          io_done,
  output wire          io_busy,
  output wire [31:0]   io_quotient,
  output wire [31:0]   io_remainder,
  input  wire          clk,
  input  wire          reset
);

  wire       [33:0]   _zz__zz_r_1;
  wire       [33:0]   _zz__zz_r_1_1;
  reg                 running;
  reg        [5:0]    counter;
  reg                 donePulse;
  reg        [32:0]   r;
  reg        [31:0]   q;
  reg        [32:0]   d;
  wire                when_UnsignedDivider_l58;
  wire       [32:0]   _zz_r;
  wire       [31:0]   _zz_q;
  wire       [33:0]   _zz_r_1;
  wire                when_UnsignedDivider_l77;
  wire                when_UnsignedDivider_l88;

  assign _zz__zz_r_1 = {1'd0, _zz_r};
  assign _zz__zz_r_1_1 = {1'd0, d};
  assign io_busy = running;
  assign io_done = donePulse;
  assign io_quotient = q;
  assign io_remainder = r[31:0];
  assign when_UnsignedDivider_l58 = (io_start && (! running));
  assign _zz_r = {r[31 : 0],q[31]};
  assign _zz_q = {q[30 : 0],1'b0};
  assign _zz_r_1 = (_zz__zz_r_1 - _zz__zz_r_1_1);
  assign when_UnsignedDivider_l77 = (! _zz_r_1[33]);
  assign when_UnsignedDivider_l88 = (counter == 6'h01);
  always @(posedge clk) begin
    if(reset) begin
      running <= 1'b0;
      counter <= 6'h0;
      donePulse <= 1'b0;
      r <= 33'h0;
      q <= 32'h0;
      d <= 33'h0;
    end else begin
      donePulse <= 1'b0;
      if(when_UnsignedDivider_l58) begin
        r <= 33'h0;
        q <= io_dividend;
        d <= {1'd0, io_divisor};
        counter <= 6'h20;
        running <= 1'b1;
      end
      if(running) begin
        if(when_UnsignedDivider_l77) begin
          r <= _zz_r_1[32:0];
          q <= (_zz_q | 32'h00000001);
        end else begin
          r <= _zz_r;
          q <= _zz_q;
        end
        counter <= (counter - 6'h01);
        if(when_UnsignedDivider_l88) begin
          running <= 1'b0;
          donePulse <= 1'b1;
        end
      end
    end
  end


endmodule

//ScratchBank_7 replaced by ScratchBank

//ScratchBank_6 replaced by ScratchBank

//ScratchBank_5 replaced by ScratchBank

//ScratchBank_4 replaced by ScratchBank

//ScratchBank_3 replaced by ScratchBank

//ScratchBank_2 replaced by ScratchBank

//ScratchBank_1 replaced by ScratchBank

module ScratchBank (
  input  wire [7:0]    io_reads_0_addr,
  input  wire          io_reads_0_en,
  output wire [31:0]   io_reads_0_data,
  input  wire [7:0]    io_reads_1_addr,
  input  wire          io_reads_1_en,
  output wire [31:0]   io_reads_1_data,
  input  wire [7:0]    io_reads_2_addr,
  input  wire          io_reads_2_en,
  output wire [31:0]   io_reads_2_data,
  input  wire [7:0]    io_write_addr,
  input  wire [31:0]   io_write_data,
  input  wire          io_write_en,
  input  wire          clk,
  input  wire          reset
);

  wire       [31:0]   replicas_0_io_rdData;
  wire       [31:0]   replicas_1_io_rdData;
  wire       [31:0]   replicas_2_io_rdData;

  BankReplica_21 replicas_0 (
    .io_rdAddr (io_reads_0_addr[7:0]      ), //i
    .io_rdEn   (io_reads_0_en             ), //i
    .io_rdData (replicas_0_io_rdData[31:0]), //o
    .io_wrAddr (io_write_addr[7:0]        ), //i
    .io_wrData (io_write_data[31:0]       ), //i
    .io_wrEn   (io_write_en               ), //i
    .clk       (clk                       ), //i
    .reset     (reset                     )  //i
  );
  BankReplica_21 replicas_1 (
    .io_rdAddr (io_reads_1_addr[7:0]      ), //i
    .io_rdEn   (io_reads_1_en             ), //i
    .io_rdData (replicas_1_io_rdData[31:0]), //o
    .io_wrAddr (io_write_addr[7:0]        ), //i
    .io_wrData (io_write_data[31:0]       ), //i
    .io_wrEn   (io_write_en               ), //i
    .clk       (clk                       ), //i
    .reset     (reset                     )  //i
  );
  BankReplica_21 replicas_2 (
    .io_rdAddr (io_reads_2_addr[7:0]      ), //i
    .io_rdEn   (io_reads_2_en             ), //i
    .io_rdData (replicas_2_io_rdData[31:0]), //o
    .io_wrAddr (io_write_addr[7:0]        ), //i
    .io_wrData (io_write_data[31:0]       ), //i
    .io_wrEn   (io_write_en               ), //i
    .clk       (clk                       ), //i
    .reset     (reset                     )  //i
  );
  assign io_reads_0_data = replicas_0_io_rdData;
  assign io_reads_1_data = replicas_1_io_rdData;
  assign io_reads_2_data = replicas_2_io_rdData;

endmodule

module StreamFifo (
  input  wire          io_push_valid,
  output wire          io_push_ready,
  input  wire [0:0]    io_push_payload,
  output reg           io_pop_valid,
  input  wire          io_pop_ready,
  output reg  [0:0]    io_pop_payload,
  input  wire          io_flush,
  output wire [2:0]    io_occupancy,
  output wire [2:0]    io_availability,
  input  wire          clk,
  input  wire          reset
);

  wire       [0:0]    logic_ram_spinal_port1;
  wire       [0:0]    _zz_logic_ram_port;
  reg                 _zz_1;
  reg                 logic_ptr_doPush;
  wire                logic_ptr_doPop;
  wire                logic_ptr_full;
  wire                logic_ptr_empty;
  reg        [2:0]    logic_ptr_push;
  reg        [2:0]    logic_ptr_pop;
  wire       [2:0]    logic_ptr_occupancy;
  wire       [2:0]    logic_ptr_popOnIo;
  wire                when_Stream_l1248;
  reg                 logic_ptr_wentUp;
  wire                io_push_fire;
  wire                logic_push_onRam_write_valid;
  wire       [1:0]    logic_push_onRam_write_payload_address;
  wire       [0:0]    logic_push_onRam_write_payload_data;
  wire                logic_pop_addressGen_valid;
  wire                logic_pop_addressGen_ready;
  wire       [1:0]    logic_pop_addressGen_payload;
  wire                logic_pop_addressGen_fire;
  wire       [0:0]    logic_pop_async_readed;
  wire                logic_pop_addressGen_translated_valid;
  wire                logic_pop_addressGen_translated_ready;
  wire       [0:0]    logic_pop_addressGen_translated_payload;
  (* ram_style = "distributed" *) reg [0:0] logic_ram [0:3];

  assign _zz_logic_ram_port = logic_push_onRam_write_payload_data;
  always @(posedge clk) begin
    if(_zz_1) begin
      logic_ram[logic_push_onRam_write_payload_address] <= _zz_logic_ram_port;
    end
  end

  assign logic_ram_spinal_port1 = logic_ram[logic_pop_addressGen_payload];
  always @(*) begin
    _zz_1 = 1'b0;
    if(logic_push_onRam_write_valid) begin
      _zz_1 = 1'b1;
    end
  end

  assign when_Stream_l1248 = (logic_ptr_doPush != logic_ptr_doPop);
  assign logic_ptr_full = (((logic_ptr_push ^ logic_ptr_popOnIo) ^ 3'b100) == 3'b000);
  assign logic_ptr_empty = (logic_ptr_push == logic_ptr_pop);
  assign logic_ptr_occupancy = (logic_ptr_push - logic_ptr_popOnIo);
  assign io_push_ready = (! logic_ptr_full);
  assign io_push_fire = (io_push_valid && io_push_ready);
  always @(*) begin
    logic_ptr_doPush = io_push_fire;
    if(logic_ptr_empty) begin
      if(io_pop_ready) begin
        logic_ptr_doPush = 1'b0;
      end
    end
  end

  assign logic_push_onRam_write_valid = io_push_fire;
  assign logic_push_onRam_write_payload_address = logic_ptr_push[1:0];
  assign logic_push_onRam_write_payload_data = io_push_payload;
  assign logic_pop_addressGen_valid = (! logic_ptr_empty);
  assign logic_pop_addressGen_payload = logic_ptr_pop[1:0];
  assign logic_pop_addressGen_fire = (logic_pop_addressGen_valid && logic_pop_addressGen_ready);
  assign logic_ptr_doPop = logic_pop_addressGen_fire;
  assign logic_pop_async_readed = logic_ram_spinal_port1;
  assign logic_pop_addressGen_translated_valid = logic_pop_addressGen_valid;
  assign logic_pop_addressGen_ready = logic_pop_addressGen_translated_ready;
  assign logic_pop_addressGen_translated_payload = logic_pop_async_readed;
  always @(*) begin
    io_pop_valid = logic_pop_addressGen_translated_valid;
    if(logic_ptr_empty) begin
      io_pop_valid = io_push_valid;
    end
  end

  assign logic_pop_addressGen_translated_ready = io_pop_ready;
  always @(*) begin
    io_pop_payload = logic_pop_addressGen_translated_payload;
    if(logic_ptr_empty) begin
      io_pop_payload = io_push_payload;
    end
  end

  assign logic_ptr_popOnIo = logic_ptr_pop;
  assign io_occupancy = logic_ptr_occupancy;
  assign io_availability = (3'b100 - logic_ptr_occupancy);
  always @(posedge clk) begin
    if(reset) begin
      logic_ptr_push <= 3'b000;
      logic_ptr_pop <= 3'b000;
      logic_ptr_wentUp <= 1'b0;
    end else begin
      if(when_Stream_l1248) begin
        logic_ptr_wentUp <= logic_ptr_doPush;
      end
      if(io_flush) begin
        logic_ptr_wentUp <= 1'b0;
      end
      if(logic_ptr_doPush) begin
        logic_ptr_push <= (logic_ptr_push + 3'b001);
      end
      if(logic_ptr_doPop) begin
        logic_ptr_pop <= (logic_ptr_pop + 3'b001);
      end
      if(io_flush) begin
        logic_ptr_push <= 3'b000;
        logic_ptr_pop <= 3'b000;
      end
    end
  end


endmodule

//BankReplica_2 replaced by BankReplica_21

//BankReplica_1 replaced by BankReplica_21

//BankReplica replaced by BankReplica_21

//BankReplica_5 replaced by BankReplica_21

//BankReplica_4 replaced by BankReplica_21

//BankReplica_3 replaced by BankReplica_21

//BankReplica_8 replaced by BankReplica_21

//BankReplica_7 replaced by BankReplica_21

//BankReplica_6 replaced by BankReplica_21

//BankReplica_11 replaced by BankReplica_21

//BankReplica_10 replaced by BankReplica_21

//BankReplica_9 replaced by BankReplica_21

//BankReplica_14 replaced by BankReplica_21

//BankReplica_13 replaced by BankReplica_21

//BankReplica_12 replaced by BankReplica_21

//BankReplica_17 replaced by BankReplica_21

//BankReplica_16 replaced by BankReplica_21

//BankReplica_15 replaced by BankReplica_21

//BankReplica_20 replaced by BankReplica_21

//BankReplica_19 replaced by BankReplica_21

//BankReplica_18 replaced by BankReplica_21

//BankReplica_23 replaced by BankReplica_21

//BankReplica_22 replaced by BankReplica_21

module BankReplica_21 (
  input  wire [7:0]    io_rdAddr,
  input  wire          io_rdEn,
  output wire [31:0]   io_rdData,
  input  wire [7:0]    io_wrAddr,
  input  wire [31:0]   io_wrData,
  input  wire          io_wrEn,
  input  wire          clk,
  input  wire          reset
);

  reg        [31:0]   mem_spinal_port0;
  wire       [31:0]   _zz_mem_port;
  reg [31:0] mem [0:191];

  assign _zz_mem_port = io_wrData;
  always @(posedge clk) begin
    if(io_rdEn) begin
      mem_spinal_port0 <= mem[io_rdAddr];
    end
    if(io_wrEn) begin
      mem[io_wrAddr] <= _zz_mem_port;
    end
  end

  assign io_rdData = mem_spinal_port0;

endmodule
