// Generator : SpinalHDL v1.10.2a    git head : a348a60b7e8b6a455c72e1536ec3d74a2ea16935
// Component : WritebackController
// Git hash  : 2b1c34e10fcfebdb7017c9a507f6d279f35a00fa

`timescale 1ns/1ps

module WritebackController (
  input  wire          io_aluWrites_0_valid,
  input  wire [10:0]   io_aluWrites_0_payload_addr,
  input  wire [31:0]   io_aluWrites_0_payload_data,
  input  wire          io_valuWrites_0_valid,
  input  wire [10:0]   io_valuWrites_0_payload_addr,
  input  wire [31:0]   io_valuWrites_0_payload_data,
  input  wire          io_valuWrites_1_valid,
  input  wire [10:0]   io_valuWrites_1_payload_addr,
  input  wire [31:0]   io_valuWrites_1_payload_data,
  input  wire          io_valuWrites_2_valid,
  input  wire [10:0]   io_valuWrites_2_payload_addr,
  input  wire [31:0]   io_valuWrites_2_payload_data,
  input  wire          io_valuWrites_3_valid,
  input  wire [10:0]   io_valuWrites_3_payload_addr,
  input  wire [31:0]   io_valuWrites_3_payload_data,
  input  wire          io_valuWrites_4_valid,
  input  wire [10:0]   io_valuWrites_4_payload_addr,
  input  wire [31:0]   io_valuWrites_4_payload_data,
  input  wire          io_valuWrites_5_valid,
  input  wire [10:0]   io_valuWrites_5_payload_addr,
  input  wire [31:0]   io_valuWrites_5_payload_data,
  input  wire          io_valuWrites_6_valid,
  input  wire [10:0]   io_valuWrites_6_payload_addr,
  input  wire [31:0]   io_valuWrites_6_payload_data,
  input  wire          io_valuWrites_7_valid,
  input  wire [10:0]   io_valuWrites_7_payload_addr,
  input  wire [31:0]   io_valuWrites_7_payload_data,
  input  wire          io_loadWrites_0_valid,
  input  wire [10:0]   io_loadWrites_0_payload_addr,
  input  wire [31:0]   io_loadWrites_0_payload_data,
  input  wire          io_constWrites_0_valid,
  input  wire [10:0]   io_constWrites_0_payload_addr,
  input  wire [31:0]   io_constWrites_0_payload_data,
  input  wire          io_vloadWrites_0_valid,
  input  wire [10:0]   io_vloadWrites_0_payload_addr,
  input  wire [31:0]   io_vloadWrites_0_payload_data,
  input  wire          io_vloadWrites_1_valid,
  input  wire [10:0]   io_vloadWrites_1_payload_addr,
  input  wire [31:0]   io_vloadWrites_1_payload_data,
  input  wire          io_vloadWrites_2_valid,
  input  wire [10:0]   io_vloadWrites_2_payload_addr,
  input  wire [31:0]   io_vloadWrites_2_payload_data,
  input  wire          io_vloadWrites_3_valid,
  input  wire [10:0]   io_vloadWrites_3_payload_addr,
  input  wire [31:0]   io_vloadWrites_3_payload_data,
  input  wire          io_vloadWrites_4_valid,
  input  wire [10:0]   io_vloadWrites_4_payload_addr,
  input  wire [31:0]   io_vloadWrites_4_payload_data,
  input  wire          io_vloadWrites_5_valid,
  input  wire [10:0]   io_vloadWrites_5_payload_addr,
  input  wire [31:0]   io_vloadWrites_5_payload_data,
  input  wire          io_vloadWrites_6_valid,
  input  wire [10:0]   io_vloadWrites_6_payload_addr,
  input  wire [31:0]   io_vloadWrites_6_payload_data,
  input  wire          io_vloadWrites_7_valid,
  input  wire [10:0]   io_vloadWrites_7_payload_addr,
  input  wire [31:0]   io_vloadWrites_7_payload_data,
  input  wire          io_flowScalarWrite_valid,
  input  wire [10:0]   io_flowScalarWrite_payload_addr,
  input  wire [31:0]   io_flowScalarWrite_payload_data,
  input  wire          io_flowVectorWrites_0_valid,
  input  wire [10:0]   io_flowVectorWrites_0_payload_addr,
  input  wire [31:0]   io_flowVectorWrites_0_payload_data,
  input  wire          io_flowVectorWrites_1_valid,
  input  wire [10:0]   io_flowVectorWrites_1_payload_addr,
  input  wire [31:0]   io_flowVectorWrites_1_payload_data,
  input  wire          io_flowVectorWrites_2_valid,
  input  wire [10:0]   io_flowVectorWrites_2_payload_addr,
  input  wire [31:0]   io_flowVectorWrites_2_payload_data,
  input  wire          io_flowVectorWrites_3_valid,
  input  wire [10:0]   io_flowVectorWrites_3_payload_addr,
  input  wire [31:0]   io_flowVectorWrites_3_payload_data,
  input  wire          io_flowVectorWrites_4_valid,
  input  wire [10:0]   io_flowVectorWrites_4_payload_addr,
  input  wire [31:0]   io_flowVectorWrites_4_payload_data,
  input  wire          io_flowVectorWrites_5_valid,
  input  wire [10:0]   io_flowVectorWrites_5_payload_addr,
  input  wire [31:0]   io_flowVectorWrites_5_payload_data,
  input  wire          io_flowVectorWrites_6_valid,
  input  wire [10:0]   io_flowVectorWrites_6_payload_addr,
  input  wire [31:0]   io_flowVectorWrites_6_payload_data,
  input  wire          io_flowVectorWrites_7_valid,
  input  wire [10:0]   io_flowVectorWrites_7_payload_addr,
  input  wire [31:0]   io_flowVectorWrites_7_payload_data,
  output wire [10:0]   io_scratchWriteAddr_0,
  output wire [10:0]   io_scratchWriteAddr_1,
  output wire [10:0]   io_scratchWriteAddr_2,
  output wire [10:0]   io_scratchWriteAddr_3,
  output wire [10:0]   io_scratchWriteAddr_4,
  output wire [10:0]   io_scratchWriteAddr_5,
  output wire [10:0]   io_scratchWriteAddr_6,
  output wire [10:0]   io_scratchWriteAddr_7,
  output wire [10:0]   io_scratchWriteAddr_8,
  output wire [10:0]   io_scratchWriteAddr_9,
  output wire [10:0]   io_scratchWriteAddr_10,
  output wire [10:0]   io_scratchWriteAddr_11,
  output wire [10:0]   io_scratchWriteAddr_12,
  output wire [10:0]   io_scratchWriteAddr_13,
  output wire [10:0]   io_scratchWriteAddr_14,
  output wire [10:0]   io_scratchWriteAddr_15,
  output wire [10:0]   io_scratchWriteAddr_16,
  output wire [10:0]   io_scratchWriteAddr_17,
  output wire [10:0]   io_scratchWriteAddr_18,
  output wire [10:0]   io_scratchWriteAddr_19,
  output wire [10:0]   io_scratchWriteAddr_20,
  output wire [10:0]   io_scratchWriteAddr_21,
  output wire [10:0]   io_scratchWriteAddr_22,
  output wire [10:0]   io_scratchWriteAddr_23,
  output wire [10:0]   io_scratchWriteAddr_24,
  output wire [10:0]   io_scratchWriteAddr_25,
  output wire [10:0]   io_scratchWriteAddr_26,
  output wire [10:0]   io_scratchWriteAddr_27,
  output wire [31:0]   io_scratchWriteData_0,
  output wire [31:0]   io_scratchWriteData_1,
  output wire [31:0]   io_scratchWriteData_2,
  output wire [31:0]   io_scratchWriteData_3,
  output wire [31:0]   io_scratchWriteData_4,
  output wire [31:0]   io_scratchWriteData_5,
  output wire [31:0]   io_scratchWriteData_6,
  output wire [31:0]   io_scratchWriteData_7,
  output wire [31:0]   io_scratchWriteData_8,
  output wire [31:0]   io_scratchWriteData_9,
  output wire [31:0]   io_scratchWriteData_10,
  output wire [31:0]   io_scratchWriteData_11,
  output wire [31:0]   io_scratchWriteData_12,
  output wire [31:0]   io_scratchWriteData_13,
  output wire [31:0]   io_scratchWriteData_14,
  output wire [31:0]   io_scratchWriteData_15,
  output wire [31:0]   io_scratchWriteData_16,
  output wire [31:0]   io_scratchWriteData_17,
  output wire [31:0]   io_scratchWriteData_18,
  output wire [31:0]   io_scratchWriteData_19,
  output wire [31:0]   io_scratchWriteData_20,
  output wire [31:0]   io_scratchWriteData_21,
  output wire [31:0]   io_scratchWriteData_22,
  output wire [31:0]   io_scratchWriteData_23,
  output wire [31:0]   io_scratchWriteData_24,
  output wire [31:0]   io_scratchWriteData_25,
  output wire [31:0]   io_scratchWriteData_26,
  output wire [31:0]   io_scratchWriteData_27,
  output wire          io_scratchWriteEn_0,
  output wire          io_scratchWriteEn_1,
  output wire          io_scratchWriteEn_2,
  output wire          io_scratchWriteEn_3,
  output wire          io_scratchWriteEn_4,
  output wire          io_scratchWriteEn_5,
  output wire          io_scratchWriteEn_6,
  output wire          io_scratchWriteEn_7,
  output wire          io_scratchWriteEn_8,
  output wire          io_scratchWriteEn_9,
  output wire          io_scratchWriteEn_10,
  output wire          io_scratchWriteEn_11,
  output wire          io_scratchWriteEn_12,
  output wire          io_scratchWriteEn_13,
  output wire          io_scratchWriteEn_14,
  output wire          io_scratchWriteEn_15,
  output wire          io_scratchWriteEn_16,
  output wire          io_scratchWriteEn_17,
  output wire          io_scratchWriteEn_18,
  output wire          io_scratchWriteEn_19,
  output wire          io_scratchWriteEn_20,
  output wire          io_scratchWriteEn_21,
  output wire          io_scratchWriteEn_22,
  output wire          io_scratchWriteEn_23,
  output wire          io_scratchWriteEn_24,
  output wire          io_scratchWriteEn_25,
  output wire          io_scratchWriteEn_26,
  output wire          io_scratchWriteEn_27,
  output reg           io_wawConflict,
  input  wire          clk,
  input  wire          reset
);

  wire                when_WritebackController_l89;
  wire                when_WritebackController_l89_1;
  wire                when_WritebackController_l89_2;
  wire                when_WritebackController_l89_3;
  wire                when_WritebackController_l89_4;
  wire                when_WritebackController_l89_5;
  wire                when_WritebackController_l89_6;
  wire                when_WritebackController_l89_7;
  wire                when_WritebackController_l89_8;
  wire                when_WritebackController_l89_9;
  wire                when_WritebackController_l89_10;
  wire                when_WritebackController_l89_11;
  wire                when_WritebackController_l89_12;
  wire                when_WritebackController_l89_13;
  wire                when_WritebackController_l89_14;
  wire                when_WritebackController_l89_15;
  wire                when_WritebackController_l89_16;
  wire                when_WritebackController_l89_17;
  wire                when_WritebackController_l89_18;
  wire                when_WritebackController_l89_19;
  wire                when_WritebackController_l89_20;
  wire                when_WritebackController_l89_21;
  wire                when_WritebackController_l89_22;
  wire                when_WritebackController_l89_23;
  wire                when_WritebackController_l89_24;
  wire                when_WritebackController_l89_25;
  wire                when_WritebackController_l89_26;
  wire                when_WritebackController_l89_27;
  wire                when_WritebackController_l89_28;
  wire                when_WritebackController_l89_29;
  wire                when_WritebackController_l89_30;
  wire                when_WritebackController_l89_31;
  wire                when_WritebackController_l89_32;
  wire                when_WritebackController_l89_33;
  wire                when_WritebackController_l89_34;
  wire                when_WritebackController_l89_35;
  wire                when_WritebackController_l89_36;
  wire                when_WritebackController_l89_37;
  wire                when_WritebackController_l89_38;
  wire                when_WritebackController_l89_39;
  wire                when_WritebackController_l89_40;
  wire                when_WritebackController_l89_41;
  wire                when_WritebackController_l89_42;
  wire                when_WritebackController_l89_43;
  wire                when_WritebackController_l89_44;
  wire                when_WritebackController_l89_45;
  wire                when_WritebackController_l89_46;
  wire                when_WritebackController_l89_47;
  wire                when_WritebackController_l89_48;
  wire                when_WritebackController_l89_49;
  wire                when_WritebackController_l89_50;
  wire                when_WritebackController_l89_51;
  wire                when_WritebackController_l89_52;
  wire                when_WritebackController_l89_53;
  wire                when_WritebackController_l89_54;
  wire                when_WritebackController_l89_55;
  wire                when_WritebackController_l89_56;
  wire                when_WritebackController_l89_57;
  wire                when_WritebackController_l89_58;
  wire                when_WritebackController_l89_59;
  wire                when_WritebackController_l89_60;
  wire                when_WritebackController_l89_61;
  wire                when_WritebackController_l89_62;
  wire                when_WritebackController_l89_63;
  wire                when_WritebackController_l89_64;
  wire                when_WritebackController_l89_65;
  wire                when_WritebackController_l89_66;
  wire                when_WritebackController_l89_67;
  wire                when_WritebackController_l89_68;
  wire                when_WritebackController_l89_69;
  wire                when_WritebackController_l89_70;
  wire                when_WritebackController_l89_71;
  wire                when_WritebackController_l89_72;
  wire                when_WritebackController_l89_73;
  wire                when_WritebackController_l89_74;
  wire                when_WritebackController_l89_75;
  wire                when_WritebackController_l89_76;
  wire                when_WritebackController_l89_77;
  wire                when_WritebackController_l89_78;
  wire                when_WritebackController_l89_79;
  wire                when_WritebackController_l89_80;
  wire                when_WritebackController_l89_81;
  wire                when_WritebackController_l89_82;
  wire                when_WritebackController_l89_83;
  wire                when_WritebackController_l89_84;
  wire                when_WritebackController_l89_85;
  wire                when_WritebackController_l89_86;
  wire                when_WritebackController_l89_87;
  wire                when_WritebackController_l89_88;
  wire                when_WritebackController_l89_89;
  wire                when_WritebackController_l89_90;
  wire                when_WritebackController_l89_91;
  wire                when_WritebackController_l89_92;
  wire                when_WritebackController_l89_93;
  wire                when_WritebackController_l89_94;
  wire                when_WritebackController_l89_95;
  wire                when_WritebackController_l89_96;
  wire                when_WritebackController_l89_97;
  wire                when_WritebackController_l89_98;
  wire                when_WritebackController_l89_99;
  wire                when_WritebackController_l89_100;
  wire                when_WritebackController_l89_101;
  wire                when_WritebackController_l89_102;
  wire                when_WritebackController_l89_103;
  wire                when_WritebackController_l89_104;
  wire                when_WritebackController_l89_105;
  wire                when_WritebackController_l89_106;
  wire                when_WritebackController_l89_107;
  wire                when_WritebackController_l89_108;
  wire                when_WritebackController_l89_109;
  wire                when_WritebackController_l89_110;
  wire                when_WritebackController_l89_111;
  wire                when_WritebackController_l89_112;
  wire                when_WritebackController_l89_113;
  wire                when_WritebackController_l89_114;
  wire                when_WritebackController_l89_115;
  wire                when_WritebackController_l89_116;
  wire                when_WritebackController_l89_117;
  wire                when_WritebackController_l89_118;
  wire                when_WritebackController_l89_119;
  wire                when_WritebackController_l89_120;
  wire                when_WritebackController_l89_121;
  wire                when_WritebackController_l89_122;
  wire                when_WritebackController_l89_123;
  wire                when_WritebackController_l89_124;
  wire                when_WritebackController_l89_125;
  wire                when_WritebackController_l89_126;
  wire                when_WritebackController_l89_127;
  wire                when_WritebackController_l89_128;
  wire                when_WritebackController_l89_129;
  wire                when_WritebackController_l89_130;
  wire                when_WritebackController_l89_131;
  wire                when_WritebackController_l89_132;
  wire                when_WritebackController_l89_133;
  wire                when_WritebackController_l89_134;
  wire                when_WritebackController_l89_135;
  wire                when_WritebackController_l89_136;
  wire                when_WritebackController_l89_137;
  wire                when_WritebackController_l89_138;
  wire                when_WritebackController_l89_139;
  wire                when_WritebackController_l89_140;
  wire                when_WritebackController_l89_141;
  wire                when_WritebackController_l89_142;
  wire                when_WritebackController_l89_143;
  wire                when_WritebackController_l89_144;
  wire                when_WritebackController_l89_145;
  wire                when_WritebackController_l89_146;
  wire                when_WritebackController_l89_147;
  wire                when_WritebackController_l89_148;
  wire                when_WritebackController_l89_149;
  wire                when_WritebackController_l89_150;
  wire                when_WritebackController_l89_151;
  wire                when_WritebackController_l89_152;
  wire                when_WritebackController_l89_153;
  wire                when_WritebackController_l89_154;
  wire                when_WritebackController_l89_155;
  wire                when_WritebackController_l89_156;
  wire                when_WritebackController_l89_157;
  wire                when_WritebackController_l89_158;
  wire                when_WritebackController_l89_159;
  wire                when_WritebackController_l89_160;
  wire                when_WritebackController_l89_161;
  wire                when_WritebackController_l89_162;
  wire                when_WritebackController_l89_163;
  wire                when_WritebackController_l89_164;
  wire                when_WritebackController_l89_165;
  wire                when_WritebackController_l89_166;
  wire                when_WritebackController_l89_167;
  wire                when_WritebackController_l89_168;
  wire                when_WritebackController_l89_169;
  wire                when_WritebackController_l89_170;
  wire                when_WritebackController_l89_171;
  wire                when_WritebackController_l89_172;
  wire                when_WritebackController_l89_173;
  wire                when_WritebackController_l89_174;
  wire                when_WritebackController_l89_175;
  wire                when_WritebackController_l89_176;
  wire                when_WritebackController_l89_177;
  wire                when_WritebackController_l89_178;
  wire                when_WritebackController_l89_179;
  wire                when_WritebackController_l89_180;
  wire                when_WritebackController_l89_181;
  wire                when_WritebackController_l89_182;
  wire                when_WritebackController_l89_183;
  wire                when_WritebackController_l89_184;
  wire                when_WritebackController_l89_185;
  wire                when_WritebackController_l89_186;
  wire                when_WritebackController_l89_187;
  wire                when_WritebackController_l89_188;
  wire                when_WritebackController_l89_189;
  wire                when_WritebackController_l89_190;
  wire                when_WritebackController_l89_191;
  wire                when_WritebackController_l89_192;
  wire                when_WritebackController_l89_193;
  wire                when_WritebackController_l89_194;
  wire                when_WritebackController_l89_195;
  wire                when_WritebackController_l89_196;
  wire                when_WritebackController_l89_197;
  wire                when_WritebackController_l89_198;
  wire                when_WritebackController_l89_199;
  wire                when_WritebackController_l89_200;
  wire                when_WritebackController_l89_201;
  wire                when_WritebackController_l89_202;
  wire                when_WritebackController_l89_203;
  wire                when_WritebackController_l89_204;
  wire                when_WritebackController_l89_205;
  wire                when_WritebackController_l89_206;
  wire                when_WritebackController_l89_207;
  wire                when_WritebackController_l89_208;
  wire                when_WritebackController_l89_209;
  wire                when_WritebackController_l89_210;
  wire                when_WritebackController_l89_211;
  wire                when_WritebackController_l89_212;
  wire                when_WritebackController_l89_213;
  wire                when_WritebackController_l89_214;
  wire                when_WritebackController_l89_215;
  wire                when_WritebackController_l89_216;
  wire                when_WritebackController_l89_217;
  wire                when_WritebackController_l89_218;
  wire                when_WritebackController_l89_219;
  wire                when_WritebackController_l89_220;
  wire                when_WritebackController_l89_221;
  wire                when_WritebackController_l89_222;
  wire                when_WritebackController_l89_223;
  wire                when_WritebackController_l89_224;
  wire                when_WritebackController_l89_225;
  wire                when_WritebackController_l89_226;
  wire                when_WritebackController_l89_227;
  wire                when_WritebackController_l89_228;
  wire                when_WritebackController_l89_229;
  wire                when_WritebackController_l89_230;
  wire                when_WritebackController_l89_231;
  wire                when_WritebackController_l89_232;
  wire                when_WritebackController_l89_233;
  wire                when_WritebackController_l89_234;
  wire                when_WritebackController_l89_235;
  wire                when_WritebackController_l89_236;
  wire                when_WritebackController_l89_237;
  wire                when_WritebackController_l89_238;
  wire                when_WritebackController_l89_239;
  wire                when_WritebackController_l89_240;
  wire                when_WritebackController_l89_241;
  wire                when_WritebackController_l89_242;
  wire                when_WritebackController_l89_243;
  wire                when_WritebackController_l89_244;
  wire                when_WritebackController_l89_245;
  wire                when_WritebackController_l89_246;
  wire                when_WritebackController_l89_247;
  wire                when_WritebackController_l89_248;
  wire                when_WritebackController_l89_249;
  wire                when_WritebackController_l89_250;
  wire                when_WritebackController_l89_251;
  wire                when_WritebackController_l89_252;
  wire                when_WritebackController_l89_253;
  wire                when_WritebackController_l89_254;
  wire                when_WritebackController_l89_255;
  wire                when_WritebackController_l89_256;
  wire                when_WritebackController_l89_257;
  wire                when_WritebackController_l89_258;
  wire                when_WritebackController_l89_259;
  wire                when_WritebackController_l89_260;
  wire                when_WritebackController_l89_261;
  wire                when_WritebackController_l89_262;
  wire                when_WritebackController_l89_263;
  wire                when_WritebackController_l89_264;
  wire                when_WritebackController_l89_265;
  wire                when_WritebackController_l89_266;
  wire                when_WritebackController_l89_267;
  wire                when_WritebackController_l89_268;
  wire                when_WritebackController_l89_269;
  wire                when_WritebackController_l89_270;
  wire                when_WritebackController_l89_271;
  wire                when_WritebackController_l89_272;
  wire                when_WritebackController_l89_273;
  wire                when_WritebackController_l89_274;
  wire                when_WritebackController_l89_275;
  wire                when_WritebackController_l89_276;
  wire                when_WritebackController_l89_277;
  wire                when_WritebackController_l89_278;
  wire                when_WritebackController_l89_279;
  wire                when_WritebackController_l89_280;
  wire                when_WritebackController_l89_281;
  wire                when_WritebackController_l89_282;
  wire                when_WritebackController_l89_283;
  wire                when_WritebackController_l89_284;
  wire                when_WritebackController_l89_285;
  wire                when_WritebackController_l89_286;
  wire                when_WritebackController_l89_287;
  wire                when_WritebackController_l89_288;
  wire                when_WritebackController_l89_289;
  wire                when_WritebackController_l89_290;
  wire                when_WritebackController_l89_291;
  wire                when_WritebackController_l89_292;
  wire                when_WritebackController_l89_293;
  wire                when_WritebackController_l89_294;
  wire                when_WritebackController_l89_295;
  wire                when_WritebackController_l89_296;
  wire                when_WritebackController_l89_297;
  wire                when_WritebackController_l89_298;
  wire                when_WritebackController_l89_299;
  wire                when_WritebackController_l89_300;
  wire                when_WritebackController_l89_301;
  wire                when_WritebackController_l89_302;
  wire                when_WritebackController_l89_303;
  wire                when_WritebackController_l89_304;
  wire                when_WritebackController_l89_305;
  wire                when_WritebackController_l89_306;
  wire                when_WritebackController_l89_307;
  wire                when_WritebackController_l89_308;
  wire                when_WritebackController_l89_309;
  wire                when_WritebackController_l89_310;
  wire                when_WritebackController_l89_311;
  wire                when_WritebackController_l89_312;
  wire                when_WritebackController_l89_313;
  wire                when_WritebackController_l89_314;
  wire                when_WritebackController_l89_315;
  wire                when_WritebackController_l89_316;
  wire                when_WritebackController_l89_317;
  wire                when_WritebackController_l89_318;
  wire                when_WritebackController_l89_319;
  wire                when_WritebackController_l89_320;
  wire                when_WritebackController_l89_321;
  wire                when_WritebackController_l89_322;
  wire                when_WritebackController_l89_323;
  wire                when_WritebackController_l89_324;
  wire                when_WritebackController_l89_325;
  wire                when_WritebackController_l89_326;
  wire                when_WritebackController_l89_327;
  wire                when_WritebackController_l89_328;
  wire                when_WritebackController_l89_329;
  wire                when_WritebackController_l89_330;
  wire                when_WritebackController_l89_331;
  wire                when_WritebackController_l89_332;
  wire                when_WritebackController_l89_333;
  wire                when_WritebackController_l89_334;
  wire                when_WritebackController_l89_335;
  wire                when_WritebackController_l89_336;
  wire                when_WritebackController_l89_337;
  wire                when_WritebackController_l89_338;
  wire                when_WritebackController_l89_339;
  wire                when_WritebackController_l89_340;
  wire                when_WritebackController_l89_341;
  wire                when_WritebackController_l89_342;
  wire                when_WritebackController_l89_343;
  wire                when_WritebackController_l89_344;
  wire                when_WritebackController_l89_345;
  wire                when_WritebackController_l89_346;
  wire                when_WritebackController_l89_347;
  wire                when_WritebackController_l89_348;
  wire                when_WritebackController_l89_349;
  wire                when_WritebackController_l89_350;
  wire                when_WritebackController_l89_351;
  wire                when_WritebackController_l89_352;
  wire                when_WritebackController_l89_353;
  wire                when_WritebackController_l89_354;
  wire                when_WritebackController_l89_355;
  wire                when_WritebackController_l89_356;
  wire                when_WritebackController_l89_357;
  wire                when_WritebackController_l89_358;
  wire                when_WritebackController_l89_359;
  wire                when_WritebackController_l89_360;
  wire                when_WritebackController_l89_361;
  wire                when_WritebackController_l89_362;
  wire                when_WritebackController_l89_363;
  wire                when_WritebackController_l89_364;
  wire                when_WritebackController_l89_365;
  wire                when_WritebackController_l89_366;
  wire                when_WritebackController_l89_367;
  wire                when_WritebackController_l89_368;
  wire                when_WritebackController_l89_369;
  wire                when_WritebackController_l89_370;
  wire                when_WritebackController_l89_371;
  wire                when_WritebackController_l89_372;
  wire                when_WritebackController_l89_373;
  wire                when_WritebackController_l89_374;
  wire                when_WritebackController_l89_375;
  wire                when_WritebackController_l89_376;
  wire                when_WritebackController_l89_377;

  assign io_scratchWriteAddr_0 = io_aluWrites_0_payload_addr;
  assign io_scratchWriteData_0 = io_aluWrites_0_payload_data;
  assign io_scratchWriteEn_0 = io_aluWrites_0_valid;
  assign io_scratchWriteAddr_1 = io_valuWrites_0_payload_addr;
  assign io_scratchWriteData_1 = io_valuWrites_0_payload_data;
  assign io_scratchWriteEn_1 = io_valuWrites_0_valid;
  assign io_scratchWriteAddr_2 = io_valuWrites_1_payload_addr;
  assign io_scratchWriteData_2 = io_valuWrites_1_payload_data;
  assign io_scratchWriteEn_2 = io_valuWrites_1_valid;
  assign io_scratchWriteAddr_3 = io_valuWrites_2_payload_addr;
  assign io_scratchWriteData_3 = io_valuWrites_2_payload_data;
  assign io_scratchWriteEn_3 = io_valuWrites_2_valid;
  assign io_scratchWriteAddr_4 = io_valuWrites_3_payload_addr;
  assign io_scratchWriteData_4 = io_valuWrites_3_payload_data;
  assign io_scratchWriteEn_4 = io_valuWrites_3_valid;
  assign io_scratchWriteAddr_5 = io_valuWrites_4_payload_addr;
  assign io_scratchWriteData_5 = io_valuWrites_4_payload_data;
  assign io_scratchWriteEn_5 = io_valuWrites_4_valid;
  assign io_scratchWriteAddr_6 = io_valuWrites_5_payload_addr;
  assign io_scratchWriteData_6 = io_valuWrites_5_payload_data;
  assign io_scratchWriteEn_6 = io_valuWrites_5_valid;
  assign io_scratchWriteAddr_7 = io_valuWrites_6_payload_addr;
  assign io_scratchWriteData_7 = io_valuWrites_6_payload_data;
  assign io_scratchWriteEn_7 = io_valuWrites_6_valid;
  assign io_scratchWriteAddr_8 = io_valuWrites_7_payload_addr;
  assign io_scratchWriteData_8 = io_valuWrites_7_payload_data;
  assign io_scratchWriteEn_8 = io_valuWrites_7_valid;
  assign io_scratchWriteAddr_9 = io_loadWrites_0_payload_addr;
  assign io_scratchWriteData_9 = io_loadWrites_0_payload_data;
  assign io_scratchWriteEn_9 = io_loadWrites_0_valid;
  assign io_scratchWriteAddr_10 = io_constWrites_0_payload_addr;
  assign io_scratchWriteData_10 = io_constWrites_0_payload_data;
  assign io_scratchWriteEn_10 = io_constWrites_0_valid;
  assign io_scratchWriteAddr_11 = io_vloadWrites_0_payload_addr;
  assign io_scratchWriteData_11 = io_vloadWrites_0_payload_data;
  assign io_scratchWriteEn_11 = io_vloadWrites_0_valid;
  assign io_scratchWriteAddr_12 = io_vloadWrites_1_payload_addr;
  assign io_scratchWriteData_12 = io_vloadWrites_1_payload_data;
  assign io_scratchWriteEn_12 = io_vloadWrites_1_valid;
  assign io_scratchWriteAddr_13 = io_vloadWrites_2_payload_addr;
  assign io_scratchWriteData_13 = io_vloadWrites_2_payload_data;
  assign io_scratchWriteEn_13 = io_vloadWrites_2_valid;
  assign io_scratchWriteAddr_14 = io_vloadWrites_3_payload_addr;
  assign io_scratchWriteData_14 = io_vloadWrites_3_payload_data;
  assign io_scratchWriteEn_14 = io_vloadWrites_3_valid;
  assign io_scratchWriteAddr_15 = io_vloadWrites_4_payload_addr;
  assign io_scratchWriteData_15 = io_vloadWrites_4_payload_data;
  assign io_scratchWriteEn_15 = io_vloadWrites_4_valid;
  assign io_scratchWriteAddr_16 = io_vloadWrites_5_payload_addr;
  assign io_scratchWriteData_16 = io_vloadWrites_5_payload_data;
  assign io_scratchWriteEn_16 = io_vloadWrites_5_valid;
  assign io_scratchWriteAddr_17 = io_vloadWrites_6_payload_addr;
  assign io_scratchWriteData_17 = io_vloadWrites_6_payload_data;
  assign io_scratchWriteEn_17 = io_vloadWrites_6_valid;
  assign io_scratchWriteAddr_18 = io_vloadWrites_7_payload_addr;
  assign io_scratchWriteData_18 = io_vloadWrites_7_payload_data;
  assign io_scratchWriteEn_18 = io_vloadWrites_7_valid;
  assign io_scratchWriteAddr_19 = io_flowScalarWrite_payload_addr;
  assign io_scratchWriteData_19 = io_flowScalarWrite_payload_data;
  assign io_scratchWriteEn_19 = io_flowScalarWrite_valid;
  assign io_scratchWriteAddr_20 = io_flowVectorWrites_0_payload_addr;
  assign io_scratchWriteData_20 = io_flowVectorWrites_0_payload_data;
  assign io_scratchWriteEn_20 = io_flowVectorWrites_0_valid;
  assign io_scratchWriteAddr_21 = io_flowVectorWrites_1_payload_addr;
  assign io_scratchWriteData_21 = io_flowVectorWrites_1_payload_data;
  assign io_scratchWriteEn_21 = io_flowVectorWrites_1_valid;
  assign io_scratchWriteAddr_22 = io_flowVectorWrites_2_payload_addr;
  assign io_scratchWriteData_22 = io_flowVectorWrites_2_payload_data;
  assign io_scratchWriteEn_22 = io_flowVectorWrites_2_valid;
  assign io_scratchWriteAddr_23 = io_flowVectorWrites_3_payload_addr;
  assign io_scratchWriteData_23 = io_flowVectorWrites_3_payload_data;
  assign io_scratchWriteEn_23 = io_flowVectorWrites_3_valid;
  assign io_scratchWriteAddr_24 = io_flowVectorWrites_4_payload_addr;
  assign io_scratchWriteData_24 = io_flowVectorWrites_4_payload_data;
  assign io_scratchWriteEn_24 = io_flowVectorWrites_4_valid;
  assign io_scratchWriteAddr_25 = io_flowVectorWrites_5_payload_addr;
  assign io_scratchWriteData_25 = io_flowVectorWrites_5_payload_data;
  assign io_scratchWriteEn_25 = io_flowVectorWrites_5_valid;
  assign io_scratchWriteAddr_26 = io_flowVectorWrites_6_payload_addr;
  assign io_scratchWriteData_26 = io_flowVectorWrites_6_payload_data;
  assign io_scratchWriteEn_26 = io_flowVectorWrites_6_valid;
  assign io_scratchWriteAddr_27 = io_flowVectorWrites_7_payload_addr;
  assign io_scratchWriteData_27 = io_flowVectorWrites_7_payload_data;
  assign io_scratchWriteEn_27 = io_flowVectorWrites_7_valid;
  always @(*) begin
    io_wawConflict = 1'b0;
    if(when_WritebackController_l89) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_1) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_2) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_3) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_4) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_5) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_6) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_7) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_8) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_9) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_10) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_11) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_12) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_13) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_14) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_15) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_16) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_17) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_18) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_19) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_20) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_21) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_22) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_23) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_24) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_25) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_26) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_27) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_28) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_29) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_30) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_31) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_32) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_33) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_34) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_35) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_36) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_37) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_38) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_39) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_40) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_41) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_42) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_43) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_44) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_45) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_46) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_47) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_48) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_49) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_50) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_51) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_52) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_53) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_54) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_55) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_56) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_57) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_58) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_59) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_60) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_61) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_62) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_63) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_64) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_65) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_66) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_67) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_68) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_69) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_70) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_71) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_72) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_73) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_74) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_75) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_76) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_77) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_78) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_79) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_80) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_81) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_82) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_83) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_84) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_85) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_86) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_87) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_88) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_89) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_90) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_91) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_92) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_93) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_94) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_95) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_96) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_97) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_98) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_99) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_100) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_101) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_102) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_103) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_104) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_105) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_106) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_107) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_108) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_109) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_110) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_111) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_112) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_113) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_114) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_115) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_116) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_117) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_118) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_119) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_120) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_121) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_122) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_123) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_124) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_125) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_126) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_127) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_128) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_129) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_130) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_131) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_132) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_133) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_134) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_135) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_136) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_137) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_138) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_139) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_140) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_141) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_142) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_143) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_144) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_145) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_146) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_147) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_148) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_149) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_150) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_151) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_152) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_153) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_154) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_155) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_156) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_157) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_158) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_159) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_160) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_161) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_162) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_163) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_164) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_165) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_166) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_167) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_168) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_169) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_170) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_171) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_172) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_173) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_174) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_175) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_176) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_177) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_178) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_179) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_180) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_181) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_182) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_183) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_184) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_185) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_186) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_187) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_188) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_189) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_190) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_191) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_192) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_193) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_194) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_195) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_196) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_197) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_198) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_199) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_200) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_201) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_202) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_203) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_204) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_205) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_206) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_207) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_208) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_209) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_210) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_211) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_212) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_213) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_214) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_215) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_216) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_217) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_218) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_219) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_220) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_221) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_222) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_223) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_224) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_225) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_226) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_227) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_228) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_229) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_230) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_231) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_232) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_233) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_234) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_235) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_236) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_237) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_238) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_239) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_240) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_241) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_242) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_243) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_244) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_245) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_246) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_247) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_248) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_249) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_250) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_251) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_252) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_253) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_254) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_255) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_256) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_257) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_258) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_259) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_260) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_261) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_262) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_263) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_264) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_265) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_266) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_267) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_268) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_269) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_270) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_271) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_272) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_273) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_274) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_275) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_276) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_277) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_278) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_279) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_280) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_281) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_282) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_283) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_284) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_285) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_286) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_287) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_288) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_289) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_290) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_291) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_292) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_293) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_294) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_295) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_296) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_297) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_298) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_299) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_300) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_301) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_302) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_303) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_304) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_305) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_306) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_307) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_308) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_309) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_310) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_311) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_312) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_313) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_314) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_315) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_316) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_317) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_318) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_319) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_320) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_321) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_322) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_323) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_324) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_325) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_326) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_327) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_328) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_329) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_330) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_331) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_332) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_333) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_334) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_335) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_336) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_337) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_338) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_339) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_340) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_341) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_342) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_343) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_344) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_345) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_346) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_347) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_348) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_349) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_350) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_351) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_352) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_353) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_354) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_355) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_356) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_357) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_358) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_359) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_360) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_361) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_362) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_363) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_364) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_365) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_366) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_367) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_368) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_369) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_370) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_371) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_372) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_373) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_374) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_375) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_376) begin
      io_wawConflict = 1'b1;
    end
    if(when_WritebackController_l89_377) begin
      io_wawConflict = 1'b1;
    end
  end

  assign when_WritebackController_l89 = ((io_aluWrites_0_valid && io_valuWrites_0_valid) && (io_aluWrites_0_payload_addr == io_valuWrites_0_payload_addr));
  assign when_WritebackController_l89_1 = ((io_aluWrites_0_valid && io_valuWrites_1_valid) && (io_aluWrites_0_payload_addr == io_valuWrites_1_payload_addr));
  assign when_WritebackController_l89_2 = ((io_aluWrites_0_valid && io_valuWrites_2_valid) && (io_aluWrites_0_payload_addr == io_valuWrites_2_payload_addr));
  assign when_WritebackController_l89_3 = ((io_aluWrites_0_valid && io_valuWrites_3_valid) && (io_aluWrites_0_payload_addr == io_valuWrites_3_payload_addr));
  assign when_WritebackController_l89_4 = ((io_aluWrites_0_valid && io_valuWrites_4_valid) && (io_aluWrites_0_payload_addr == io_valuWrites_4_payload_addr));
  assign when_WritebackController_l89_5 = ((io_aluWrites_0_valid && io_valuWrites_5_valid) && (io_aluWrites_0_payload_addr == io_valuWrites_5_payload_addr));
  assign when_WritebackController_l89_6 = ((io_aluWrites_0_valid && io_valuWrites_6_valid) && (io_aluWrites_0_payload_addr == io_valuWrites_6_payload_addr));
  assign when_WritebackController_l89_7 = ((io_aluWrites_0_valid && io_valuWrites_7_valid) && (io_aluWrites_0_payload_addr == io_valuWrites_7_payload_addr));
  assign when_WritebackController_l89_8 = ((io_aluWrites_0_valid && io_loadWrites_0_valid) && (io_aluWrites_0_payload_addr == io_loadWrites_0_payload_addr));
  assign when_WritebackController_l89_9 = ((io_aluWrites_0_valid && io_constWrites_0_valid) && (io_aluWrites_0_payload_addr == io_constWrites_0_payload_addr));
  assign when_WritebackController_l89_10 = ((io_aluWrites_0_valid && io_vloadWrites_0_valid) && (io_aluWrites_0_payload_addr == io_vloadWrites_0_payload_addr));
  assign when_WritebackController_l89_11 = ((io_aluWrites_0_valid && io_vloadWrites_1_valid) && (io_aluWrites_0_payload_addr == io_vloadWrites_1_payload_addr));
  assign when_WritebackController_l89_12 = ((io_aluWrites_0_valid && io_vloadWrites_2_valid) && (io_aluWrites_0_payload_addr == io_vloadWrites_2_payload_addr));
  assign when_WritebackController_l89_13 = ((io_aluWrites_0_valid && io_vloadWrites_3_valid) && (io_aluWrites_0_payload_addr == io_vloadWrites_3_payload_addr));
  assign when_WritebackController_l89_14 = ((io_aluWrites_0_valid && io_vloadWrites_4_valid) && (io_aluWrites_0_payload_addr == io_vloadWrites_4_payload_addr));
  assign when_WritebackController_l89_15 = ((io_aluWrites_0_valid && io_vloadWrites_5_valid) && (io_aluWrites_0_payload_addr == io_vloadWrites_5_payload_addr));
  assign when_WritebackController_l89_16 = ((io_aluWrites_0_valid && io_vloadWrites_6_valid) && (io_aluWrites_0_payload_addr == io_vloadWrites_6_payload_addr));
  assign when_WritebackController_l89_17 = ((io_aluWrites_0_valid && io_vloadWrites_7_valid) && (io_aluWrites_0_payload_addr == io_vloadWrites_7_payload_addr));
  assign when_WritebackController_l89_18 = ((io_aluWrites_0_valid && io_flowScalarWrite_valid) && (io_aluWrites_0_payload_addr == io_flowScalarWrite_payload_addr));
  assign when_WritebackController_l89_19 = ((io_aluWrites_0_valid && io_flowVectorWrites_0_valid) && (io_aluWrites_0_payload_addr == io_flowVectorWrites_0_payload_addr));
  assign when_WritebackController_l89_20 = ((io_aluWrites_0_valid && io_flowVectorWrites_1_valid) && (io_aluWrites_0_payload_addr == io_flowVectorWrites_1_payload_addr));
  assign when_WritebackController_l89_21 = ((io_aluWrites_0_valid && io_flowVectorWrites_2_valid) && (io_aluWrites_0_payload_addr == io_flowVectorWrites_2_payload_addr));
  assign when_WritebackController_l89_22 = ((io_aluWrites_0_valid && io_flowVectorWrites_3_valid) && (io_aluWrites_0_payload_addr == io_flowVectorWrites_3_payload_addr));
  assign when_WritebackController_l89_23 = ((io_aluWrites_0_valid && io_flowVectorWrites_4_valid) && (io_aluWrites_0_payload_addr == io_flowVectorWrites_4_payload_addr));
  assign when_WritebackController_l89_24 = ((io_aluWrites_0_valid && io_flowVectorWrites_5_valid) && (io_aluWrites_0_payload_addr == io_flowVectorWrites_5_payload_addr));
  assign when_WritebackController_l89_25 = ((io_aluWrites_0_valid && io_flowVectorWrites_6_valid) && (io_aluWrites_0_payload_addr == io_flowVectorWrites_6_payload_addr));
  assign when_WritebackController_l89_26 = ((io_aluWrites_0_valid && io_flowVectorWrites_7_valid) && (io_aluWrites_0_payload_addr == io_flowVectorWrites_7_payload_addr));
  assign when_WritebackController_l89_27 = ((io_valuWrites_0_valid && io_valuWrites_1_valid) && (io_valuWrites_0_payload_addr == io_valuWrites_1_payload_addr));
  assign when_WritebackController_l89_28 = ((io_valuWrites_0_valid && io_valuWrites_2_valid) && (io_valuWrites_0_payload_addr == io_valuWrites_2_payload_addr));
  assign when_WritebackController_l89_29 = ((io_valuWrites_0_valid && io_valuWrites_3_valid) && (io_valuWrites_0_payload_addr == io_valuWrites_3_payload_addr));
  assign when_WritebackController_l89_30 = ((io_valuWrites_0_valid && io_valuWrites_4_valid) && (io_valuWrites_0_payload_addr == io_valuWrites_4_payload_addr));
  assign when_WritebackController_l89_31 = ((io_valuWrites_0_valid && io_valuWrites_5_valid) && (io_valuWrites_0_payload_addr == io_valuWrites_5_payload_addr));
  assign when_WritebackController_l89_32 = ((io_valuWrites_0_valid && io_valuWrites_6_valid) && (io_valuWrites_0_payload_addr == io_valuWrites_6_payload_addr));
  assign when_WritebackController_l89_33 = ((io_valuWrites_0_valid && io_valuWrites_7_valid) && (io_valuWrites_0_payload_addr == io_valuWrites_7_payload_addr));
  assign when_WritebackController_l89_34 = ((io_valuWrites_0_valid && io_loadWrites_0_valid) && (io_valuWrites_0_payload_addr == io_loadWrites_0_payload_addr));
  assign when_WritebackController_l89_35 = ((io_valuWrites_0_valid && io_constWrites_0_valid) && (io_valuWrites_0_payload_addr == io_constWrites_0_payload_addr));
  assign when_WritebackController_l89_36 = ((io_valuWrites_0_valid && io_vloadWrites_0_valid) && (io_valuWrites_0_payload_addr == io_vloadWrites_0_payload_addr));
  assign when_WritebackController_l89_37 = ((io_valuWrites_0_valid && io_vloadWrites_1_valid) && (io_valuWrites_0_payload_addr == io_vloadWrites_1_payload_addr));
  assign when_WritebackController_l89_38 = ((io_valuWrites_0_valid && io_vloadWrites_2_valid) && (io_valuWrites_0_payload_addr == io_vloadWrites_2_payload_addr));
  assign when_WritebackController_l89_39 = ((io_valuWrites_0_valid && io_vloadWrites_3_valid) && (io_valuWrites_0_payload_addr == io_vloadWrites_3_payload_addr));
  assign when_WritebackController_l89_40 = ((io_valuWrites_0_valid && io_vloadWrites_4_valid) && (io_valuWrites_0_payload_addr == io_vloadWrites_4_payload_addr));
  assign when_WritebackController_l89_41 = ((io_valuWrites_0_valid && io_vloadWrites_5_valid) && (io_valuWrites_0_payload_addr == io_vloadWrites_5_payload_addr));
  assign when_WritebackController_l89_42 = ((io_valuWrites_0_valid && io_vloadWrites_6_valid) && (io_valuWrites_0_payload_addr == io_vloadWrites_6_payload_addr));
  assign when_WritebackController_l89_43 = ((io_valuWrites_0_valid && io_vloadWrites_7_valid) && (io_valuWrites_0_payload_addr == io_vloadWrites_7_payload_addr));
  assign when_WritebackController_l89_44 = ((io_valuWrites_0_valid && io_flowScalarWrite_valid) && (io_valuWrites_0_payload_addr == io_flowScalarWrite_payload_addr));
  assign when_WritebackController_l89_45 = ((io_valuWrites_0_valid && io_flowVectorWrites_0_valid) && (io_valuWrites_0_payload_addr == io_flowVectorWrites_0_payload_addr));
  assign when_WritebackController_l89_46 = ((io_valuWrites_0_valid && io_flowVectorWrites_1_valid) && (io_valuWrites_0_payload_addr == io_flowVectorWrites_1_payload_addr));
  assign when_WritebackController_l89_47 = ((io_valuWrites_0_valid && io_flowVectorWrites_2_valid) && (io_valuWrites_0_payload_addr == io_flowVectorWrites_2_payload_addr));
  assign when_WritebackController_l89_48 = ((io_valuWrites_0_valid && io_flowVectorWrites_3_valid) && (io_valuWrites_0_payload_addr == io_flowVectorWrites_3_payload_addr));
  assign when_WritebackController_l89_49 = ((io_valuWrites_0_valid && io_flowVectorWrites_4_valid) && (io_valuWrites_0_payload_addr == io_flowVectorWrites_4_payload_addr));
  assign when_WritebackController_l89_50 = ((io_valuWrites_0_valid && io_flowVectorWrites_5_valid) && (io_valuWrites_0_payload_addr == io_flowVectorWrites_5_payload_addr));
  assign when_WritebackController_l89_51 = ((io_valuWrites_0_valid && io_flowVectorWrites_6_valid) && (io_valuWrites_0_payload_addr == io_flowVectorWrites_6_payload_addr));
  assign when_WritebackController_l89_52 = ((io_valuWrites_0_valid && io_flowVectorWrites_7_valid) && (io_valuWrites_0_payload_addr == io_flowVectorWrites_7_payload_addr));
  assign when_WritebackController_l89_53 = ((io_valuWrites_1_valid && io_valuWrites_2_valid) && (io_valuWrites_1_payload_addr == io_valuWrites_2_payload_addr));
  assign when_WritebackController_l89_54 = ((io_valuWrites_1_valid && io_valuWrites_3_valid) && (io_valuWrites_1_payload_addr == io_valuWrites_3_payload_addr));
  assign when_WritebackController_l89_55 = ((io_valuWrites_1_valid && io_valuWrites_4_valid) && (io_valuWrites_1_payload_addr == io_valuWrites_4_payload_addr));
  assign when_WritebackController_l89_56 = ((io_valuWrites_1_valid && io_valuWrites_5_valid) && (io_valuWrites_1_payload_addr == io_valuWrites_5_payload_addr));
  assign when_WritebackController_l89_57 = ((io_valuWrites_1_valid && io_valuWrites_6_valid) && (io_valuWrites_1_payload_addr == io_valuWrites_6_payload_addr));
  assign when_WritebackController_l89_58 = ((io_valuWrites_1_valid && io_valuWrites_7_valid) && (io_valuWrites_1_payload_addr == io_valuWrites_7_payload_addr));
  assign when_WritebackController_l89_59 = ((io_valuWrites_1_valid && io_loadWrites_0_valid) && (io_valuWrites_1_payload_addr == io_loadWrites_0_payload_addr));
  assign when_WritebackController_l89_60 = ((io_valuWrites_1_valid && io_constWrites_0_valid) && (io_valuWrites_1_payload_addr == io_constWrites_0_payload_addr));
  assign when_WritebackController_l89_61 = ((io_valuWrites_1_valid && io_vloadWrites_0_valid) && (io_valuWrites_1_payload_addr == io_vloadWrites_0_payload_addr));
  assign when_WritebackController_l89_62 = ((io_valuWrites_1_valid && io_vloadWrites_1_valid) && (io_valuWrites_1_payload_addr == io_vloadWrites_1_payload_addr));
  assign when_WritebackController_l89_63 = ((io_valuWrites_1_valid && io_vloadWrites_2_valid) && (io_valuWrites_1_payload_addr == io_vloadWrites_2_payload_addr));
  assign when_WritebackController_l89_64 = ((io_valuWrites_1_valid && io_vloadWrites_3_valid) && (io_valuWrites_1_payload_addr == io_vloadWrites_3_payload_addr));
  assign when_WritebackController_l89_65 = ((io_valuWrites_1_valid && io_vloadWrites_4_valid) && (io_valuWrites_1_payload_addr == io_vloadWrites_4_payload_addr));
  assign when_WritebackController_l89_66 = ((io_valuWrites_1_valid && io_vloadWrites_5_valid) && (io_valuWrites_1_payload_addr == io_vloadWrites_5_payload_addr));
  assign when_WritebackController_l89_67 = ((io_valuWrites_1_valid && io_vloadWrites_6_valid) && (io_valuWrites_1_payload_addr == io_vloadWrites_6_payload_addr));
  assign when_WritebackController_l89_68 = ((io_valuWrites_1_valid && io_vloadWrites_7_valid) && (io_valuWrites_1_payload_addr == io_vloadWrites_7_payload_addr));
  assign when_WritebackController_l89_69 = ((io_valuWrites_1_valid && io_flowScalarWrite_valid) && (io_valuWrites_1_payload_addr == io_flowScalarWrite_payload_addr));
  assign when_WritebackController_l89_70 = ((io_valuWrites_1_valid && io_flowVectorWrites_0_valid) && (io_valuWrites_1_payload_addr == io_flowVectorWrites_0_payload_addr));
  assign when_WritebackController_l89_71 = ((io_valuWrites_1_valid && io_flowVectorWrites_1_valid) && (io_valuWrites_1_payload_addr == io_flowVectorWrites_1_payload_addr));
  assign when_WritebackController_l89_72 = ((io_valuWrites_1_valid && io_flowVectorWrites_2_valid) && (io_valuWrites_1_payload_addr == io_flowVectorWrites_2_payload_addr));
  assign when_WritebackController_l89_73 = ((io_valuWrites_1_valid && io_flowVectorWrites_3_valid) && (io_valuWrites_1_payload_addr == io_flowVectorWrites_3_payload_addr));
  assign when_WritebackController_l89_74 = ((io_valuWrites_1_valid && io_flowVectorWrites_4_valid) && (io_valuWrites_1_payload_addr == io_flowVectorWrites_4_payload_addr));
  assign when_WritebackController_l89_75 = ((io_valuWrites_1_valid && io_flowVectorWrites_5_valid) && (io_valuWrites_1_payload_addr == io_flowVectorWrites_5_payload_addr));
  assign when_WritebackController_l89_76 = ((io_valuWrites_1_valid && io_flowVectorWrites_6_valid) && (io_valuWrites_1_payload_addr == io_flowVectorWrites_6_payload_addr));
  assign when_WritebackController_l89_77 = ((io_valuWrites_1_valid && io_flowVectorWrites_7_valid) && (io_valuWrites_1_payload_addr == io_flowVectorWrites_7_payload_addr));
  assign when_WritebackController_l89_78 = ((io_valuWrites_2_valid && io_valuWrites_3_valid) && (io_valuWrites_2_payload_addr == io_valuWrites_3_payload_addr));
  assign when_WritebackController_l89_79 = ((io_valuWrites_2_valid && io_valuWrites_4_valid) && (io_valuWrites_2_payload_addr == io_valuWrites_4_payload_addr));
  assign when_WritebackController_l89_80 = ((io_valuWrites_2_valid && io_valuWrites_5_valid) && (io_valuWrites_2_payload_addr == io_valuWrites_5_payload_addr));
  assign when_WritebackController_l89_81 = ((io_valuWrites_2_valid && io_valuWrites_6_valid) && (io_valuWrites_2_payload_addr == io_valuWrites_6_payload_addr));
  assign when_WritebackController_l89_82 = ((io_valuWrites_2_valid && io_valuWrites_7_valid) && (io_valuWrites_2_payload_addr == io_valuWrites_7_payload_addr));
  assign when_WritebackController_l89_83 = ((io_valuWrites_2_valid && io_loadWrites_0_valid) && (io_valuWrites_2_payload_addr == io_loadWrites_0_payload_addr));
  assign when_WritebackController_l89_84 = ((io_valuWrites_2_valid && io_constWrites_0_valid) && (io_valuWrites_2_payload_addr == io_constWrites_0_payload_addr));
  assign when_WritebackController_l89_85 = ((io_valuWrites_2_valid && io_vloadWrites_0_valid) && (io_valuWrites_2_payload_addr == io_vloadWrites_0_payload_addr));
  assign when_WritebackController_l89_86 = ((io_valuWrites_2_valid && io_vloadWrites_1_valid) && (io_valuWrites_2_payload_addr == io_vloadWrites_1_payload_addr));
  assign when_WritebackController_l89_87 = ((io_valuWrites_2_valid && io_vloadWrites_2_valid) && (io_valuWrites_2_payload_addr == io_vloadWrites_2_payload_addr));
  assign when_WritebackController_l89_88 = ((io_valuWrites_2_valid && io_vloadWrites_3_valid) && (io_valuWrites_2_payload_addr == io_vloadWrites_3_payload_addr));
  assign when_WritebackController_l89_89 = ((io_valuWrites_2_valid && io_vloadWrites_4_valid) && (io_valuWrites_2_payload_addr == io_vloadWrites_4_payload_addr));
  assign when_WritebackController_l89_90 = ((io_valuWrites_2_valid && io_vloadWrites_5_valid) && (io_valuWrites_2_payload_addr == io_vloadWrites_5_payload_addr));
  assign when_WritebackController_l89_91 = ((io_valuWrites_2_valid && io_vloadWrites_6_valid) && (io_valuWrites_2_payload_addr == io_vloadWrites_6_payload_addr));
  assign when_WritebackController_l89_92 = ((io_valuWrites_2_valid && io_vloadWrites_7_valid) && (io_valuWrites_2_payload_addr == io_vloadWrites_7_payload_addr));
  assign when_WritebackController_l89_93 = ((io_valuWrites_2_valid && io_flowScalarWrite_valid) && (io_valuWrites_2_payload_addr == io_flowScalarWrite_payload_addr));
  assign when_WritebackController_l89_94 = ((io_valuWrites_2_valid && io_flowVectorWrites_0_valid) && (io_valuWrites_2_payload_addr == io_flowVectorWrites_0_payload_addr));
  assign when_WritebackController_l89_95 = ((io_valuWrites_2_valid && io_flowVectorWrites_1_valid) && (io_valuWrites_2_payload_addr == io_flowVectorWrites_1_payload_addr));
  assign when_WritebackController_l89_96 = ((io_valuWrites_2_valid && io_flowVectorWrites_2_valid) && (io_valuWrites_2_payload_addr == io_flowVectorWrites_2_payload_addr));
  assign when_WritebackController_l89_97 = ((io_valuWrites_2_valid && io_flowVectorWrites_3_valid) && (io_valuWrites_2_payload_addr == io_flowVectorWrites_3_payload_addr));
  assign when_WritebackController_l89_98 = ((io_valuWrites_2_valid && io_flowVectorWrites_4_valid) && (io_valuWrites_2_payload_addr == io_flowVectorWrites_4_payload_addr));
  assign when_WritebackController_l89_99 = ((io_valuWrites_2_valid && io_flowVectorWrites_5_valid) && (io_valuWrites_2_payload_addr == io_flowVectorWrites_5_payload_addr));
  assign when_WritebackController_l89_100 = ((io_valuWrites_2_valid && io_flowVectorWrites_6_valid) && (io_valuWrites_2_payload_addr == io_flowVectorWrites_6_payload_addr));
  assign when_WritebackController_l89_101 = ((io_valuWrites_2_valid && io_flowVectorWrites_7_valid) && (io_valuWrites_2_payload_addr == io_flowVectorWrites_7_payload_addr));
  assign when_WritebackController_l89_102 = ((io_valuWrites_3_valid && io_valuWrites_4_valid) && (io_valuWrites_3_payload_addr == io_valuWrites_4_payload_addr));
  assign when_WritebackController_l89_103 = ((io_valuWrites_3_valid && io_valuWrites_5_valid) && (io_valuWrites_3_payload_addr == io_valuWrites_5_payload_addr));
  assign when_WritebackController_l89_104 = ((io_valuWrites_3_valid && io_valuWrites_6_valid) && (io_valuWrites_3_payload_addr == io_valuWrites_6_payload_addr));
  assign when_WritebackController_l89_105 = ((io_valuWrites_3_valid && io_valuWrites_7_valid) && (io_valuWrites_3_payload_addr == io_valuWrites_7_payload_addr));
  assign when_WritebackController_l89_106 = ((io_valuWrites_3_valid && io_loadWrites_0_valid) && (io_valuWrites_3_payload_addr == io_loadWrites_0_payload_addr));
  assign when_WritebackController_l89_107 = ((io_valuWrites_3_valid && io_constWrites_0_valid) && (io_valuWrites_3_payload_addr == io_constWrites_0_payload_addr));
  assign when_WritebackController_l89_108 = ((io_valuWrites_3_valid && io_vloadWrites_0_valid) && (io_valuWrites_3_payload_addr == io_vloadWrites_0_payload_addr));
  assign when_WritebackController_l89_109 = ((io_valuWrites_3_valid && io_vloadWrites_1_valid) && (io_valuWrites_3_payload_addr == io_vloadWrites_1_payload_addr));
  assign when_WritebackController_l89_110 = ((io_valuWrites_3_valid && io_vloadWrites_2_valid) && (io_valuWrites_3_payload_addr == io_vloadWrites_2_payload_addr));
  assign when_WritebackController_l89_111 = ((io_valuWrites_3_valid && io_vloadWrites_3_valid) && (io_valuWrites_3_payload_addr == io_vloadWrites_3_payload_addr));
  assign when_WritebackController_l89_112 = ((io_valuWrites_3_valid && io_vloadWrites_4_valid) && (io_valuWrites_3_payload_addr == io_vloadWrites_4_payload_addr));
  assign when_WritebackController_l89_113 = ((io_valuWrites_3_valid && io_vloadWrites_5_valid) && (io_valuWrites_3_payload_addr == io_vloadWrites_5_payload_addr));
  assign when_WritebackController_l89_114 = ((io_valuWrites_3_valid && io_vloadWrites_6_valid) && (io_valuWrites_3_payload_addr == io_vloadWrites_6_payload_addr));
  assign when_WritebackController_l89_115 = ((io_valuWrites_3_valid && io_vloadWrites_7_valid) && (io_valuWrites_3_payload_addr == io_vloadWrites_7_payload_addr));
  assign when_WritebackController_l89_116 = ((io_valuWrites_3_valid && io_flowScalarWrite_valid) && (io_valuWrites_3_payload_addr == io_flowScalarWrite_payload_addr));
  assign when_WritebackController_l89_117 = ((io_valuWrites_3_valid && io_flowVectorWrites_0_valid) && (io_valuWrites_3_payload_addr == io_flowVectorWrites_0_payload_addr));
  assign when_WritebackController_l89_118 = ((io_valuWrites_3_valid && io_flowVectorWrites_1_valid) && (io_valuWrites_3_payload_addr == io_flowVectorWrites_1_payload_addr));
  assign when_WritebackController_l89_119 = ((io_valuWrites_3_valid && io_flowVectorWrites_2_valid) && (io_valuWrites_3_payload_addr == io_flowVectorWrites_2_payload_addr));
  assign when_WritebackController_l89_120 = ((io_valuWrites_3_valid && io_flowVectorWrites_3_valid) && (io_valuWrites_3_payload_addr == io_flowVectorWrites_3_payload_addr));
  assign when_WritebackController_l89_121 = ((io_valuWrites_3_valid && io_flowVectorWrites_4_valid) && (io_valuWrites_3_payload_addr == io_flowVectorWrites_4_payload_addr));
  assign when_WritebackController_l89_122 = ((io_valuWrites_3_valid && io_flowVectorWrites_5_valid) && (io_valuWrites_3_payload_addr == io_flowVectorWrites_5_payload_addr));
  assign when_WritebackController_l89_123 = ((io_valuWrites_3_valid && io_flowVectorWrites_6_valid) && (io_valuWrites_3_payload_addr == io_flowVectorWrites_6_payload_addr));
  assign when_WritebackController_l89_124 = ((io_valuWrites_3_valid && io_flowVectorWrites_7_valid) && (io_valuWrites_3_payload_addr == io_flowVectorWrites_7_payload_addr));
  assign when_WritebackController_l89_125 = ((io_valuWrites_4_valid && io_valuWrites_5_valid) && (io_valuWrites_4_payload_addr == io_valuWrites_5_payload_addr));
  assign when_WritebackController_l89_126 = ((io_valuWrites_4_valid && io_valuWrites_6_valid) && (io_valuWrites_4_payload_addr == io_valuWrites_6_payload_addr));
  assign when_WritebackController_l89_127 = ((io_valuWrites_4_valid && io_valuWrites_7_valid) && (io_valuWrites_4_payload_addr == io_valuWrites_7_payload_addr));
  assign when_WritebackController_l89_128 = ((io_valuWrites_4_valid && io_loadWrites_0_valid) && (io_valuWrites_4_payload_addr == io_loadWrites_0_payload_addr));
  assign when_WritebackController_l89_129 = ((io_valuWrites_4_valid && io_constWrites_0_valid) && (io_valuWrites_4_payload_addr == io_constWrites_0_payload_addr));
  assign when_WritebackController_l89_130 = ((io_valuWrites_4_valid && io_vloadWrites_0_valid) && (io_valuWrites_4_payload_addr == io_vloadWrites_0_payload_addr));
  assign when_WritebackController_l89_131 = ((io_valuWrites_4_valid && io_vloadWrites_1_valid) && (io_valuWrites_4_payload_addr == io_vloadWrites_1_payload_addr));
  assign when_WritebackController_l89_132 = ((io_valuWrites_4_valid && io_vloadWrites_2_valid) && (io_valuWrites_4_payload_addr == io_vloadWrites_2_payload_addr));
  assign when_WritebackController_l89_133 = ((io_valuWrites_4_valid && io_vloadWrites_3_valid) && (io_valuWrites_4_payload_addr == io_vloadWrites_3_payload_addr));
  assign when_WritebackController_l89_134 = ((io_valuWrites_4_valid && io_vloadWrites_4_valid) && (io_valuWrites_4_payload_addr == io_vloadWrites_4_payload_addr));
  assign when_WritebackController_l89_135 = ((io_valuWrites_4_valid && io_vloadWrites_5_valid) && (io_valuWrites_4_payload_addr == io_vloadWrites_5_payload_addr));
  assign when_WritebackController_l89_136 = ((io_valuWrites_4_valid && io_vloadWrites_6_valid) && (io_valuWrites_4_payload_addr == io_vloadWrites_6_payload_addr));
  assign when_WritebackController_l89_137 = ((io_valuWrites_4_valid && io_vloadWrites_7_valid) && (io_valuWrites_4_payload_addr == io_vloadWrites_7_payload_addr));
  assign when_WritebackController_l89_138 = ((io_valuWrites_4_valid && io_flowScalarWrite_valid) && (io_valuWrites_4_payload_addr == io_flowScalarWrite_payload_addr));
  assign when_WritebackController_l89_139 = ((io_valuWrites_4_valid && io_flowVectorWrites_0_valid) && (io_valuWrites_4_payload_addr == io_flowVectorWrites_0_payload_addr));
  assign when_WritebackController_l89_140 = ((io_valuWrites_4_valid && io_flowVectorWrites_1_valid) && (io_valuWrites_4_payload_addr == io_flowVectorWrites_1_payload_addr));
  assign when_WritebackController_l89_141 = ((io_valuWrites_4_valid && io_flowVectorWrites_2_valid) && (io_valuWrites_4_payload_addr == io_flowVectorWrites_2_payload_addr));
  assign when_WritebackController_l89_142 = ((io_valuWrites_4_valid && io_flowVectorWrites_3_valid) && (io_valuWrites_4_payload_addr == io_flowVectorWrites_3_payload_addr));
  assign when_WritebackController_l89_143 = ((io_valuWrites_4_valid && io_flowVectorWrites_4_valid) && (io_valuWrites_4_payload_addr == io_flowVectorWrites_4_payload_addr));
  assign when_WritebackController_l89_144 = ((io_valuWrites_4_valid && io_flowVectorWrites_5_valid) && (io_valuWrites_4_payload_addr == io_flowVectorWrites_5_payload_addr));
  assign when_WritebackController_l89_145 = ((io_valuWrites_4_valid && io_flowVectorWrites_6_valid) && (io_valuWrites_4_payload_addr == io_flowVectorWrites_6_payload_addr));
  assign when_WritebackController_l89_146 = ((io_valuWrites_4_valid && io_flowVectorWrites_7_valid) && (io_valuWrites_4_payload_addr == io_flowVectorWrites_7_payload_addr));
  assign when_WritebackController_l89_147 = ((io_valuWrites_5_valid && io_valuWrites_6_valid) && (io_valuWrites_5_payload_addr == io_valuWrites_6_payload_addr));
  assign when_WritebackController_l89_148 = ((io_valuWrites_5_valid && io_valuWrites_7_valid) && (io_valuWrites_5_payload_addr == io_valuWrites_7_payload_addr));
  assign when_WritebackController_l89_149 = ((io_valuWrites_5_valid && io_loadWrites_0_valid) && (io_valuWrites_5_payload_addr == io_loadWrites_0_payload_addr));
  assign when_WritebackController_l89_150 = ((io_valuWrites_5_valid && io_constWrites_0_valid) && (io_valuWrites_5_payload_addr == io_constWrites_0_payload_addr));
  assign when_WritebackController_l89_151 = ((io_valuWrites_5_valid && io_vloadWrites_0_valid) && (io_valuWrites_5_payload_addr == io_vloadWrites_0_payload_addr));
  assign when_WritebackController_l89_152 = ((io_valuWrites_5_valid && io_vloadWrites_1_valid) && (io_valuWrites_5_payload_addr == io_vloadWrites_1_payload_addr));
  assign when_WritebackController_l89_153 = ((io_valuWrites_5_valid && io_vloadWrites_2_valid) && (io_valuWrites_5_payload_addr == io_vloadWrites_2_payload_addr));
  assign when_WritebackController_l89_154 = ((io_valuWrites_5_valid && io_vloadWrites_3_valid) && (io_valuWrites_5_payload_addr == io_vloadWrites_3_payload_addr));
  assign when_WritebackController_l89_155 = ((io_valuWrites_5_valid && io_vloadWrites_4_valid) && (io_valuWrites_5_payload_addr == io_vloadWrites_4_payload_addr));
  assign when_WritebackController_l89_156 = ((io_valuWrites_5_valid && io_vloadWrites_5_valid) && (io_valuWrites_5_payload_addr == io_vloadWrites_5_payload_addr));
  assign when_WritebackController_l89_157 = ((io_valuWrites_5_valid && io_vloadWrites_6_valid) && (io_valuWrites_5_payload_addr == io_vloadWrites_6_payload_addr));
  assign when_WritebackController_l89_158 = ((io_valuWrites_5_valid && io_vloadWrites_7_valid) && (io_valuWrites_5_payload_addr == io_vloadWrites_7_payload_addr));
  assign when_WritebackController_l89_159 = ((io_valuWrites_5_valid && io_flowScalarWrite_valid) && (io_valuWrites_5_payload_addr == io_flowScalarWrite_payload_addr));
  assign when_WritebackController_l89_160 = ((io_valuWrites_5_valid && io_flowVectorWrites_0_valid) && (io_valuWrites_5_payload_addr == io_flowVectorWrites_0_payload_addr));
  assign when_WritebackController_l89_161 = ((io_valuWrites_5_valid && io_flowVectorWrites_1_valid) && (io_valuWrites_5_payload_addr == io_flowVectorWrites_1_payload_addr));
  assign when_WritebackController_l89_162 = ((io_valuWrites_5_valid && io_flowVectorWrites_2_valid) && (io_valuWrites_5_payload_addr == io_flowVectorWrites_2_payload_addr));
  assign when_WritebackController_l89_163 = ((io_valuWrites_5_valid && io_flowVectorWrites_3_valid) && (io_valuWrites_5_payload_addr == io_flowVectorWrites_3_payload_addr));
  assign when_WritebackController_l89_164 = ((io_valuWrites_5_valid && io_flowVectorWrites_4_valid) && (io_valuWrites_5_payload_addr == io_flowVectorWrites_4_payload_addr));
  assign when_WritebackController_l89_165 = ((io_valuWrites_5_valid && io_flowVectorWrites_5_valid) && (io_valuWrites_5_payload_addr == io_flowVectorWrites_5_payload_addr));
  assign when_WritebackController_l89_166 = ((io_valuWrites_5_valid && io_flowVectorWrites_6_valid) && (io_valuWrites_5_payload_addr == io_flowVectorWrites_6_payload_addr));
  assign when_WritebackController_l89_167 = ((io_valuWrites_5_valid && io_flowVectorWrites_7_valid) && (io_valuWrites_5_payload_addr == io_flowVectorWrites_7_payload_addr));
  assign when_WritebackController_l89_168 = ((io_valuWrites_6_valid && io_valuWrites_7_valid) && (io_valuWrites_6_payload_addr == io_valuWrites_7_payload_addr));
  assign when_WritebackController_l89_169 = ((io_valuWrites_6_valid && io_loadWrites_0_valid) && (io_valuWrites_6_payload_addr == io_loadWrites_0_payload_addr));
  assign when_WritebackController_l89_170 = ((io_valuWrites_6_valid && io_constWrites_0_valid) && (io_valuWrites_6_payload_addr == io_constWrites_0_payload_addr));
  assign when_WritebackController_l89_171 = ((io_valuWrites_6_valid && io_vloadWrites_0_valid) && (io_valuWrites_6_payload_addr == io_vloadWrites_0_payload_addr));
  assign when_WritebackController_l89_172 = ((io_valuWrites_6_valid && io_vloadWrites_1_valid) && (io_valuWrites_6_payload_addr == io_vloadWrites_1_payload_addr));
  assign when_WritebackController_l89_173 = ((io_valuWrites_6_valid && io_vloadWrites_2_valid) && (io_valuWrites_6_payload_addr == io_vloadWrites_2_payload_addr));
  assign when_WritebackController_l89_174 = ((io_valuWrites_6_valid && io_vloadWrites_3_valid) && (io_valuWrites_6_payload_addr == io_vloadWrites_3_payload_addr));
  assign when_WritebackController_l89_175 = ((io_valuWrites_6_valid && io_vloadWrites_4_valid) && (io_valuWrites_6_payload_addr == io_vloadWrites_4_payload_addr));
  assign when_WritebackController_l89_176 = ((io_valuWrites_6_valid && io_vloadWrites_5_valid) && (io_valuWrites_6_payload_addr == io_vloadWrites_5_payload_addr));
  assign when_WritebackController_l89_177 = ((io_valuWrites_6_valid && io_vloadWrites_6_valid) && (io_valuWrites_6_payload_addr == io_vloadWrites_6_payload_addr));
  assign when_WritebackController_l89_178 = ((io_valuWrites_6_valid && io_vloadWrites_7_valid) && (io_valuWrites_6_payload_addr == io_vloadWrites_7_payload_addr));
  assign when_WritebackController_l89_179 = ((io_valuWrites_6_valid && io_flowScalarWrite_valid) && (io_valuWrites_6_payload_addr == io_flowScalarWrite_payload_addr));
  assign when_WritebackController_l89_180 = ((io_valuWrites_6_valid && io_flowVectorWrites_0_valid) && (io_valuWrites_6_payload_addr == io_flowVectorWrites_0_payload_addr));
  assign when_WritebackController_l89_181 = ((io_valuWrites_6_valid && io_flowVectorWrites_1_valid) && (io_valuWrites_6_payload_addr == io_flowVectorWrites_1_payload_addr));
  assign when_WritebackController_l89_182 = ((io_valuWrites_6_valid && io_flowVectorWrites_2_valid) && (io_valuWrites_6_payload_addr == io_flowVectorWrites_2_payload_addr));
  assign when_WritebackController_l89_183 = ((io_valuWrites_6_valid && io_flowVectorWrites_3_valid) && (io_valuWrites_6_payload_addr == io_flowVectorWrites_3_payload_addr));
  assign when_WritebackController_l89_184 = ((io_valuWrites_6_valid && io_flowVectorWrites_4_valid) && (io_valuWrites_6_payload_addr == io_flowVectorWrites_4_payload_addr));
  assign when_WritebackController_l89_185 = ((io_valuWrites_6_valid && io_flowVectorWrites_5_valid) && (io_valuWrites_6_payload_addr == io_flowVectorWrites_5_payload_addr));
  assign when_WritebackController_l89_186 = ((io_valuWrites_6_valid && io_flowVectorWrites_6_valid) && (io_valuWrites_6_payload_addr == io_flowVectorWrites_6_payload_addr));
  assign when_WritebackController_l89_187 = ((io_valuWrites_6_valid && io_flowVectorWrites_7_valid) && (io_valuWrites_6_payload_addr == io_flowVectorWrites_7_payload_addr));
  assign when_WritebackController_l89_188 = ((io_valuWrites_7_valid && io_loadWrites_0_valid) && (io_valuWrites_7_payload_addr == io_loadWrites_0_payload_addr));
  assign when_WritebackController_l89_189 = ((io_valuWrites_7_valid && io_constWrites_0_valid) && (io_valuWrites_7_payload_addr == io_constWrites_0_payload_addr));
  assign when_WritebackController_l89_190 = ((io_valuWrites_7_valid && io_vloadWrites_0_valid) && (io_valuWrites_7_payload_addr == io_vloadWrites_0_payload_addr));
  assign when_WritebackController_l89_191 = ((io_valuWrites_7_valid && io_vloadWrites_1_valid) && (io_valuWrites_7_payload_addr == io_vloadWrites_1_payload_addr));
  assign when_WritebackController_l89_192 = ((io_valuWrites_7_valid && io_vloadWrites_2_valid) && (io_valuWrites_7_payload_addr == io_vloadWrites_2_payload_addr));
  assign when_WritebackController_l89_193 = ((io_valuWrites_7_valid && io_vloadWrites_3_valid) && (io_valuWrites_7_payload_addr == io_vloadWrites_3_payload_addr));
  assign when_WritebackController_l89_194 = ((io_valuWrites_7_valid && io_vloadWrites_4_valid) && (io_valuWrites_7_payload_addr == io_vloadWrites_4_payload_addr));
  assign when_WritebackController_l89_195 = ((io_valuWrites_7_valid && io_vloadWrites_5_valid) && (io_valuWrites_7_payload_addr == io_vloadWrites_5_payload_addr));
  assign when_WritebackController_l89_196 = ((io_valuWrites_7_valid && io_vloadWrites_6_valid) && (io_valuWrites_7_payload_addr == io_vloadWrites_6_payload_addr));
  assign when_WritebackController_l89_197 = ((io_valuWrites_7_valid && io_vloadWrites_7_valid) && (io_valuWrites_7_payload_addr == io_vloadWrites_7_payload_addr));
  assign when_WritebackController_l89_198 = ((io_valuWrites_7_valid && io_flowScalarWrite_valid) && (io_valuWrites_7_payload_addr == io_flowScalarWrite_payload_addr));
  assign when_WritebackController_l89_199 = ((io_valuWrites_7_valid && io_flowVectorWrites_0_valid) && (io_valuWrites_7_payload_addr == io_flowVectorWrites_0_payload_addr));
  assign when_WritebackController_l89_200 = ((io_valuWrites_7_valid && io_flowVectorWrites_1_valid) && (io_valuWrites_7_payload_addr == io_flowVectorWrites_1_payload_addr));
  assign when_WritebackController_l89_201 = ((io_valuWrites_7_valid && io_flowVectorWrites_2_valid) && (io_valuWrites_7_payload_addr == io_flowVectorWrites_2_payload_addr));
  assign when_WritebackController_l89_202 = ((io_valuWrites_7_valid && io_flowVectorWrites_3_valid) && (io_valuWrites_7_payload_addr == io_flowVectorWrites_3_payload_addr));
  assign when_WritebackController_l89_203 = ((io_valuWrites_7_valid && io_flowVectorWrites_4_valid) && (io_valuWrites_7_payload_addr == io_flowVectorWrites_4_payload_addr));
  assign when_WritebackController_l89_204 = ((io_valuWrites_7_valid && io_flowVectorWrites_5_valid) && (io_valuWrites_7_payload_addr == io_flowVectorWrites_5_payload_addr));
  assign when_WritebackController_l89_205 = ((io_valuWrites_7_valid && io_flowVectorWrites_6_valid) && (io_valuWrites_7_payload_addr == io_flowVectorWrites_6_payload_addr));
  assign when_WritebackController_l89_206 = ((io_valuWrites_7_valid && io_flowVectorWrites_7_valid) && (io_valuWrites_7_payload_addr == io_flowVectorWrites_7_payload_addr));
  assign when_WritebackController_l89_207 = ((io_loadWrites_0_valid && io_constWrites_0_valid) && (io_loadWrites_0_payload_addr == io_constWrites_0_payload_addr));
  assign when_WritebackController_l89_208 = ((io_loadWrites_0_valid && io_vloadWrites_0_valid) && (io_loadWrites_0_payload_addr == io_vloadWrites_0_payload_addr));
  assign when_WritebackController_l89_209 = ((io_loadWrites_0_valid && io_vloadWrites_1_valid) && (io_loadWrites_0_payload_addr == io_vloadWrites_1_payload_addr));
  assign when_WritebackController_l89_210 = ((io_loadWrites_0_valid && io_vloadWrites_2_valid) && (io_loadWrites_0_payload_addr == io_vloadWrites_2_payload_addr));
  assign when_WritebackController_l89_211 = ((io_loadWrites_0_valid && io_vloadWrites_3_valid) && (io_loadWrites_0_payload_addr == io_vloadWrites_3_payload_addr));
  assign when_WritebackController_l89_212 = ((io_loadWrites_0_valid && io_vloadWrites_4_valid) && (io_loadWrites_0_payload_addr == io_vloadWrites_4_payload_addr));
  assign when_WritebackController_l89_213 = ((io_loadWrites_0_valid && io_vloadWrites_5_valid) && (io_loadWrites_0_payload_addr == io_vloadWrites_5_payload_addr));
  assign when_WritebackController_l89_214 = ((io_loadWrites_0_valid && io_vloadWrites_6_valid) && (io_loadWrites_0_payload_addr == io_vloadWrites_6_payload_addr));
  assign when_WritebackController_l89_215 = ((io_loadWrites_0_valid && io_vloadWrites_7_valid) && (io_loadWrites_0_payload_addr == io_vloadWrites_7_payload_addr));
  assign when_WritebackController_l89_216 = ((io_loadWrites_0_valid && io_flowScalarWrite_valid) && (io_loadWrites_0_payload_addr == io_flowScalarWrite_payload_addr));
  assign when_WritebackController_l89_217 = ((io_loadWrites_0_valid && io_flowVectorWrites_0_valid) && (io_loadWrites_0_payload_addr == io_flowVectorWrites_0_payload_addr));
  assign when_WritebackController_l89_218 = ((io_loadWrites_0_valid && io_flowVectorWrites_1_valid) && (io_loadWrites_0_payload_addr == io_flowVectorWrites_1_payload_addr));
  assign when_WritebackController_l89_219 = ((io_loadWrites_0_valid && io_flowVectorWrites_2_valid) && (io_loadWrites_0_payload_addr == io_flowVectorWrites_2_payload_addr));
  assign when_WritebackController_l89_220 = ((io_loadWrites_0_valid && io_flowVectorWrites_3_valid) && (io_loadWrites_0_payload_addr == io_flowVectorWrites_3_payload_addr));
  assign when_WritebackController_l89_221 = ((io_loadWrites_0_valid && io_flowVectorWrites_4_valid) && (io_loadWrites_0_payload_addr == io_flowVectorWrites_4_payload_addr));
  assign when_WritebackController_l89_222 = ((io_loadWrites_0_valid && io_flowVectorWrites_5_valid) && (io_loadWrites_0_payload_addr == io_flowVectorWrites_5_payload_addr));
  assign when_WritebackController_l89_223 = ((io_loadWrites_0_valid && io_flowVectorWrites_6_valid) && (io_loadWrites_0_payload_addr == io_flowVectorWrites_6_payload_addr));
  assign when_WritebackController_l89_224 = ((io_loadWrites_0_valid && io_flowVectorWrites_7_valid) && (io_loadWrites_0_payload_addr == io_flowVectorWrites_7_payload_addr));
  assign when_WritebackController_l89_225 = ((io_constWrites_0_valid && io_vloadWrites_0_valid) && (io_constWrites_0_payload_addr == io_vloadWrites_0_payload_addr));
  assign when_WritebackController_l89_226 = ((io_constWrites_0_valid && io_vloadWrites_1_valid) && (io_constWrites_0_payload_addr == io_vloadWrites_1_payload_addr));
  assign when_WritebackController_l89_227 = ((io_constWrites_0_valid && io_vloadWrites_2_valid) && (io_constWrites_0_payload_addr == io_vloadWrites_2_payload_addr));
  assign when_WritebackController_l89_228 = ((io_constWrites_0_valid && io_vloadWrites_3_valid) && (io_constWrites_0_payload_addr == io_vloadWrites_3_payload_addr));
  assign when_WritebackController_l89_229 = ((io_constWrites_0_valid && io_vloadWrites_4_valid) && (io_constWrites_0_payload_addr == io_vloadWrites_4_payload_addr));
  assign when_WritebackController_l89_230 = ((io_constWrites_0_valid && io_vloadWrites_5_valid) && (io_constWrites_0_payload_addr == io_vloadWrites_5_payload_addr));
  assign when_WritebackController_l89_231 = ((io_constWrites_0_valid && io_vloadWrites_6_valid) && (io_constWrites_0_payload_addr == io_vloadWrites_6_payload_addr));
  assign when_WritebackController_l89_232 = ((io_constWrites_0_valid && io_vloadWrites_7_valid) && (io_constWrites_0_payload_addr == io_vloadWrites_7_payload_addr));
  assign when_WritebackController_l89_233 = ((io_constWrites_0_valid && io_flowScalarWrite_valid) && (io_constWrites_0_payload_addr == io_flowScalarWrite_payload_addr));
  assign when_WritebackController_l89_234 = ((io_constWrites_0_valid && io_flowVectorWrites_0_valid) && (io_constWrites_0_payload_addr == io_flowVectorWrites_0_payload_addr));
  assign when_WritebackController_l89_235 = ((io_constWrites_0_valid && io_flowVectorWrites_1_valid) && (io_constWrites_0_payload_addr == io_flowVectorWrites_1_payload_addr));
  assign when_WritebackController_l89_236 = ((io_constWrites_0_valid && io_flowVectorWrites_2_valid) && (io_constWrites_0_payload_addr == io_flowVectorWrites_2_payload_addr));
  assign when_WritebackController_l89_237 = ((io_constWrites_0_valid && io_flowVectorWrites_3_valid) && (io_constWrites_0_payload_addr == io_flowVectorWrites_3_payload_addr));
  assign when_WritebackController_l89_238 = ((io_constWrites_0_valid && io_flowVectorWrites_4_valid) && (io_constWrites_0_payload_addr == io_flowVectorWrites_4_payload_addr));
  assign when_WritebackController_l89_239 = ((io_constWrites_0_valid && io_flowVectorWrites_5_valid) && (io_constWrites_0_payload_addr == io_flowVectorWrites_5_payload_addr));
  assign when_WritebackController_l89_240 = ((io_constWrites_0_valid && io_flowVectorWrites_6_valid) && (io_constWrites_0_payload_addr == io_flowVectorWrites_6_payload_addr));
  assign when_WritebackController_l89_241 = ((io_constWrites_0_valid && io_flowVectorWrites_7_valid) && (io_constWrites_0_payload_addr == io_flowVectorWrites_7_payload_addr));
  assign when_WritebackController_l89_242 = ((io_vloadWrites_0_valid && io_vloadWrites_1_valid) && (io_vloadWrites_0_payload_addr == io_vloadWrites_1_payload_addr));
  assign when_WritebackController_l89_243 = ((io_vloadWrites_0_valid && io_vloadWrites_2_valid) && (io_vloadWrites_0_payload_addr == io_vloadWrites_2_payload_addr));
  assign when_WritebackController_l89_244 = ((io_vloadWrites_0_valid && io_vloadWrites_3_valid) && (io_vloadWrites_0_payload_addr == io_vloadWrites_3_payload_addr));
  assign when_WritebackController_l89_245 = ((io_vloadWrites_0_valid && io_vloadWrites_4_valid) && (io_vloadWrites_0_payload_addr == io_vloadWrites_4_payload_addr));
  assign when_WritebackController_l89_246 = ((io_vloadWrites_0_valid && io_vloadWrites_5_valid) && (io_vloadWrites_0_payload_addr == io_vloadWrites_5_payload_addr));
  assign when_WritebackController_l89_247 = ((io_vloadWrites_0_valid && io_vloadWrites_6_valid) && (io_vloadWrites_0_payload_addr == io_vloadWrites_6_payload_addr));
  assign when_WritebackController_l89_248 = ((io_vloadWrites_0_valid && io_vloadWrites_7_valid) && (io_vloadWrites_0_payload_addr == io_vloadWrites_7_payload_addr));
  assign when_WritebackController_l89_249 = ((io_vloadWrites_0_valid && io_flowScalarWrite_valid) && (io_vloadWrites_0_payload_addr == io_flowScalarWrite_payload_addr));
  assign when_WritebackController_l89_250 = ((io_vloadWrites_0_valid && io_flowVectorWrites_0_valid) && (io_vloadWrites_0_payload_addr == io_flowVectorWrites_0_payload_addr));
  assign when_WritebackController_l89_251 = ((io_vloadWrites_0_valid && io_flowVectorWrites_1_valid) && (io_vloadWrites_0_payload_addr == io_flowVectorWrites_1_payload_addr));
  assign when_WritebackController_l89_252 = ((io_vloadWrites_0_valid && io_flowVectorWrites_2_valid) && (io_vloadWrites_0_payload_addr == io_flowVectorWrites_2_payload_addr));
  assign when_WritebackController_l89_253 = ((io_vloadWrites_0_valid && io_flowVectorWrites_3_valid) && (io_vloadWrites_0_payload_addr == io_flowVectorWrites_3_payload_addr));
  assign when_WritebackController_l89_254 = ((io_vloadWrites_0_valid && io_flowVectorWrites_4_valid) && (io_vloadWrites_0_payload_addr == io_flowVectorWrites_4_payload_addr));
  assign when_WritebackController_l89_255 = ((io_vloadWrites_0_valid && io_flowVectorWrites_5_valid) && (io_vloadWrites_0_payload_addr == io_flowVectorWrites_5_payload_addr));
  assign when_WritebackController_l89_256 = ((io_vloadWrites_0_valid && io_flowVectorWrites_6_valid) && (io_vloadWrites_0_payload_addr == io_flowVectorWrites_6_payload_addr));
  assign when_WritebackController_l89_257 = ((io_vloadWrites_0_valid && io_flowVectorWrites_7_valid) && (io_vloadWrites_0_payload_addr == io_flowVectorWrites_7_payload_addr));
  assign when_WritebackController_l89_258 = ((io_vloadWrites_1_valid && io_vloadWrites_2_valid) && (io_vloadWrites_1_payload_addr == io_vloadWrites_2_payload_addr));
  assign when_WritebackController_l89_259 = ((io_vloadWrites_1_valid && io_vloadWrites_3_valid) && (io_vloadWrites_1_payload_addr == io_vloadWrites_3_payload_addr));
  assign when_WritebackController_l89_260 = ((io_vloadWrites_1_valid && io_vloadWrites_4_valid) && (io_vloadWrites_1_payload_addr == io_vloadWrites_4_payload_addr));
  assign when_WritebackController_l89_261 = ((io_vloadWrites_1_valid && io_vloadWrites_5_valid) && (io_vloadWrites_1_payload_addr == io_vloadWrites_5_payload_addr));
  assign when_WritebackController_l89_262 = ((io_vloadWrites_1_valid && io_vloadWrites_6_valid) && (io_vloadWrites_1_payload_addr == io_vloadWrites_6_payload_addr));
  assign when_WritebackController_l89_263 = ((io_vloadWrites_1_valid && io_vloadWrites_7_valid) && (io_vloadWrites_1_payload_addr == io_vloadWrites_7_payload_addr));
  assign when_WritebackController_l89_264 = ((io_vloadWrites_1_valid && io_flowScalarWrite_valid) && (io_vloadWrites_1_payload_addr == io_flowScalarWrite_payload_addr));
  assign when_WritebackController_l89_265 = ((io_vloadWrites_1_valid && io_flowVectorWrites_0_valid) && (io_vloadWrites_1_payload_addr == io_flowVectorWrites_0_payload_addr));
  assign when_WritebackController_l89_266 = ((io_vloadWrites_1_valid && io_flowVectorWrites_1_valid) && (io_vloadWrites_1_payload_addr == io_flowVectorWrites_1_payload_addr));
  assign when_WritebackController_l89_267 = ((io_vloadWrites_1_valid && io_flowVectorWrites_2_valid) && (io_vloadWrites_1_payload_addr == io_flowVectorWrites_2_payload_addr));
  assign when_WritebackController_l89_268 = ((io_vloadWrites_1_valid && io_flowVectorWrites_3_valid) && (io_vloadWrites_1_payload_addr == io_flowVectorWrites_3_payload_addr));
  assign when_WritebackController_l89_269 = ((io_vloadWrites_1_valid && io_flowVectorWrites_4_valid) && (io_vloadWrites_1_payload_addr == io_flowVectorWrites_4_payload_addr));
  assign when_WritebackController_l89_270 = ((io_vloadWrites_1_valid && io_flowVectorWrites_5_valid) && (io_vloadWrites_1_payload_addr == io_flowVectorWrites_5_payload_addr));
  assign when_WritebackController_l89_271 = ((io_vloadWrites_1_valid && io_flowVectorWrites_6_valid) && (io_vloadWrites_1_payload_addr == io_flowVectorWrites_6_payload_addr));
  assign when_WritebackController_l89_272 = ((io_vloadWrites_1_valid && io_flowVectorWrites_7_valid) && (io_vloadWrites_1_payload_addr == io_flowVectorWrites_7_payload_addr));
  assign when_WritebackController_l89_273 = ((io_vloadWrites_2_valid && io_vloadWrites_3_valid) && (io_vloadWrites_2_payload_addr == io_vloadWrites_3_payload_addr));
  assign when_WritebackController_l89_274 = ((io_vloadWrites_2_valid && io_vloadWrites_4_valid) && (io_vloadWrites_2_payload_addr == io_vloadWrites_4_payload_addr));
  assign when_WritebackController_l89_275 = ((io_vloadWrites_2_valid && io_vloadWrites_5_valid) && (io_vloadWrites_2_payload_addr == io_vloadWrites_5_payload_addr));
  assign when_WritebackController_l89_276 = ((io_vloadWrites_2_valid && io_vloadWrites_6_valid) && (io_vloadWrites_2_payload_addr == io_vloadWrites_6_payload_addr));
  assign when_WritebackController_l89_277 = ((io_vloadWrites_2_valid && io_vloadWrites_7_valid) && (io_vloadWrites_2_payload_addr == io_vloadWrites_7_payload_addr));
  assign when_WritebackController_l89_278 = ((io_vloadWrites_2_valid && io_flowScalarWrite_valid) && (io_vloadWrites_2_payload_addr == io_flowScalarWrite_payload_addr));
  assign when_WritebackController_l89_279 = ((io_vloadWrites_2_valid && io_flowVectorWrites_0_valid) && (io_vloadWrites_2_payload_addr == io_flowVectorWrites_0_payload_addr));
  assign when_WritebackController_l89_280 = ((io_vloadWrites_2_valid && io_flowVectorWrites_1_valid) && (io_vloadWrites_2_payload_addr == io_flowVectorWrites_1_payload_addr));
  assign when_WritebackController_l89_281 = ((io_vloadWrites_2_valid && io_flowVectorWrites_2_valid) && (io_vloadWrites_2_payload_addr == io_flowVectorWrites_2_payload_addr));
  assign when_WritebackController_l89_282 = ((io_vloadWrites_2_valid && io_flowVectorWrites_3_valid) && (io_vloadWrites_2_payload_addr == io_flowVectorWrites_3_payload_addr));
  assign when_WritebackController_l89_283 = ((io_vloadWrites_2_valid && io_flowVectorWrites_4_valid) && (io_vloadWrites_2_payload_addr == io_flowVectorWrites_4_payload_addr));
  assign when_WritebackController_l89_284 = ((io_vloadWrites_2_valid && io_flowVectorWrites_5_valid) && (io_vloadWrites_2_payload_addr == io_flowVectorWrites_5_payload_addr));
  assign when_WritebackController_l89_285 = ((io_vloadWrites_2_valid && io_flowVectorWrites_6_valid) && (io_vloadWrites_2_payload_addr == io_flowVectorWrites_6_payload_addr));
  assign when_WritebackController_l89_286 = ((io_vloadWrites_2_valid && io_flowVectorWrites_7_valid) && (io_vloadWrites_2_payload_addr == io_flowVectorWrites_7_payload_addr));
  assign when_WritebackController_l89_287 = ((io_vloadWrites_3_valid && io_vloadWrites_4_valid) && (io_vloadWrites_3_payload_addr == io_vloadWrites_4_payload_addr));
  assign when_WritebackController_l89_288 = ((io_vloadWrites_3_valid && io_vloadWrites_5_valid) && (io_vloadWrites_3_payload_addr == io_vloadWrites_5_payload_addr));
  assign when_WritebackController_l89_289 = ((io_vloadWrites_3_valid && io_vloadWrites_6_valid) && (io_vloadWrites_3_payload_addr == io_vloadWrites_6_payload_addr));
  assign when_WritebackController_l89_290 = ((io_vloadWrites_3_valid && io_vloadWrites_7_valid) && (io_vloadWrites_3_payload_addr == io_vloadWrites_7_payload_addr));
  assign when_WritebackController_l89_291 = ((io_vloadWrites_3_valid && io_flowScalarWrite_valid) && (io_vloadWrites_3_payload_addr == io_flowScalarWrite_payload_addr));
  assign when_WritebackController_l89_292 = ((io_vloadWrites_3_valid && io_flowVectorWrites_0_valid) && (io_vloadWrites_3_payload_addr == io_flowVectorWrites_0_payload_addr));
  assign when_WritebackController_l89_293 = ((io_vloadWrites_3_valid && io_flowVectorWrites_1_valid) && (io_vloadWrites_3_payload_addr == io_flowVectorWrites_1_payload_addr));
  assign when_WritebackController_l89_294 = ((io_vloadWrites_3_valid && io_flowVectorWrites_2_valid) && (io_vloadWrites_3_payload_addr == io_flowVectorWrites_2_payload_addr));
  assign when_WritebackController_l89_295 = ((io_vloadWrites_3_valid && io_flowVectorWrites_3_valid) && (io_vloadWrites_3_payload_addr == io_flowVectorWrites_3_payload_addr));
  assign when_WritebackController_l89_296 = ((io_vloadWrites_3_valid && io_flowVectorWrites_4_valid) && (io_vloadWrites_3_payload_addr == io_flowVectorWrites_4_payload_addr));
  assign when_WritebackController_l89_297 = ((io_vloadWrites_3_valid && io_flowVectorWrites_5_valid) && (io_vloadWrites_3_payload_addr == io_flowVectorWrites_5_payload_addr));
  assign when_WritebackController_l89_298 = ((io_vloadWrites_3_valid && io_flowVectorWrites_6_valid) && (io_vloadWrites_3_payload_addr == io_flowVectorWrites_6_payload_addr));
  assign when_WritebackController_l89_299 = ((io_vloadWrites_3_valid && io_flowVectorWrites_7_valid) && (io_vloadWrites_3_payload_addr == io_flowVectorWrites_7_payload_addr));
  assign when_WritebackController_l89_300 = ((io_vloadWrites_4_valid && io_vloadWrites_5_valid) && (io_vloadWrites_4_payload_addr == io_vloadWrites_5_payload_addr));
  assign when_WritebackController_l89_301 = ((io_vloadWrites_4_valid && io_vloadWrites_6_valid) && (io_vloadWrites_4_payload_addr == io_vloadWrites_6_payload_addr));
  assign when_WritebackController_l89_302 = ((io_vloadWrites_4_valid && io_vloadWrites_7_valid) && (io_vloadWrites_4_payload_addr == io_vloadWrites_7_payload_addr));
  assign when_WritebackController_l89_303 = ((io_vloadWrites_4_valid && io_flowScalarWrite_valid) && (io_vloadWrites_4_payload_addr == io_flowScalarWrite_payload_addr));
  assign when_WritebackController_l89_304 = ((io_vloadWrites_4_valid && io_flowVectorWrites_0_valid) && (io_vloadWrites_4_payload_addr == io_flowVectorWrites_0_payload_addr));
  assign when_WritebackController_l89_305 = ((io_vloadWrites_4_valid && io_flowVectorWrites_1_valid) && (io_vloadWrites_4_payload_addr == io_flowVectorWrites_1_payload_addr));
  assign when_WritebackController_l89_306 = ((io_vloadWrites_4_valid && io_flowVectorWrites_2_valid) && (io_vloadWrites_4_payload_addr == io_flowVectorWrites_2_payload_addr));
  assign when_WritebackController_l89_307 = ((io_vloadWrites_4_valid && io_flowVectorWrites_3_valid) && (io_vloadWrites_4_payload_addr == io_flowVectorWrites_3_payload_addr));
  assign when_WritebackController_l89_308 = ((io_vloadWrites_4_valid && io_flowVectorWrites_4_valid) && (io_vloadWrites_4_payload_addr == io_flowVectorWrites_4_payload_addr));
  assign when_WritebackController_l89_309 = ((io_vloadWrites_4_valid && io_flowVectorWrites_5_valid) && (io_vloadWrites_4_payload_addr == io_flowVectorWrites_5_payload_addr));
  assign when_WritebackController_l89_310 = ((io_vloadWrites_4_valid && io_flowVectorWrites_6_valid) && (io_vloadWrites_4_payload_addr == io_flowVectorWrites_6_payload_addr));
  assign when_WritebackController_l89_311 = ((io_vloadWrites_4_valid && io_flowVectorWrites_7_valid) && (io_vloadWrites_4_payload_addr == io_flowVectorWrites_7_payload_addr));
  assign when_WritebackController_l89_312 = ((io_vloadWrites_5_valid && io_vloadWrites_6_valid) && (io_vloadWrites_5_payload_addr == io_vloadWrites_6_payload_addr));
  assign when_WritebackController_l89_313 = ((io_vloadWrites_5_valid && io_vloadWrites_7_valid) && (io_vloadWrites_5_payload_addr == io_vloadWrites_7_payload_addr));
  assign when_WritebackController_l89_314 = ((io_vloadWrites_5_valid && io_flowScalarWrite_valid) && (io_vloadWrites_5_payload_addr == io_flowScalarWrite_payload_addr));
  assign when_WritebackController_l89_315 = ((io_vloadWrites_5_valid && io_flowVectorWrites_0_valid) && (io_vloadWrites_5_payload_addr == io_flowVectorWrites_0_payload_addr));
  assign when_WritebackController_l89_316 = ((io_vloadWrites_5_valid && io_flowVectorWrites_1_valid) && (io_vloadWrites_5_payload_addr == io_flowVectorWrites_1_payload_addr));
  assign when_WritebackController_l89_317 = ((io_vloadWrites_5_valid && io_flowVectorWrites_2_valid) && (io_vloadWrites_5_payload_addr == io_flowVectorWrites_2_payload_addr));
  assign when_WritebackController_l89_318 = ((io_vloadWrites_5_valid && io_flowVectorWrites_3_valid) && (io_vloadWrites_5_payload_addr == io_flowVectorWrites_3_payload_addr));
  assign when_WritebackController_l89_319 = ((io_vloadWrites_5_valid && io_flowVectorWrites_4_valid) && (io_vloadWrites_5_payload_addr == io_flowVectorWrites_4_payload_addr));
  assign when_WritebackController_l89_320 = ((io_vloadWrites_5_valid && io_flowVectorWrites_5_valid) && (io_vloadWrites_5_payload_addr == io_flowVectorWrites_5_payload_addr));
  assign when_WritebackController_l89_321 = ((io_vloadWrites_5_valid && io_flowVectorWrites_6_valid) && (io_vloadWrites_5_payload_addr == io_flowVectorWrites_6_payload_addr));
  assign when_WritebackController_l89_322 = ((io_vloadWrites_5_valid && io_flowVectorWrites_7_valid) && (io_vloadWrites_5_payload_addr == io_flowVectorWrites_7_payload_addr));
  assign when_WritebackController_l89_323 = ((io_vloadWrites_6_valid && io_vloadWrites_7_valid) && (io_vloadWrites_6_payload_addr == io_vloadWrites_7_payload_addr));
  assign when_WritebackController_l89_324 = ((io_vloadWrites_6_valid && io_flowScalarWrite_valid) && (io_vloadWrites_6_payload_addr == io_flowScalarWrite_payload_addr));
  assign when_WritebackController_l89_325 = ((io_vloadWrites_6_valid && io_flowVectorWrites_0_valid) && (io_vloadWrites_6_payload_addr == io_flowVectorWrites_0_payload_addr));
  assign when_WritebackController_l89_326 = ((io_vloadWrites_6_valid && io_flowVectorWrites_1_valid) && (io_vloadWrites_6_payload_addr == io_flowVectorWrites_1_payload_addr));
  assign when_WritebackController_l89_327 = ((io_vloadWrites_6_valid && io_flowVectorWrites_2_valid) && (io_vloadWrites_6_payload_addr == io_flowVectorWrites_2_payload_addr));
  assign when_WritebackController_l89_328 = ((io_vloadWrites_6_valid && io_flowVectorWrites_3_valid) && (io_vloadWrites_6_payload_addr == io_flowVectorWrites_3_payload_addr));
  assign when_WritebackController_l89_329 = ((io_vloadWrites_6_valid && io_flowVectorWrites_4_valid) && (io_vloadWrites_6_payload_addr == io_flowVectorWrites_4_payload_addr));
  assign when_WritebackController_l89_330 = ((io_vloadWrites_6_valid && io_flowVectorWrites_5_valid) && (io_vloadWrites_6_payload_addr == io_flowVectorWrites_5_payload_addr));
  assign when_WritebackController_l89_331 = ((io_vloadWrites_6_valid && io_flowVectorWrites_6_valid) && (io_vloadWrites_6_payload_addr == io_flowVectorWrites_6_payload_addr));
  assign when_WritebackController_l89_332 = ((io_vloadWrites_6_valid && io_flowVectorWrites_7_valid) && (io_vloadWrites_6_payload_addr == io_flowVectorWrites_7_payload_addr));
  assign when_WritebackController_l89_333 = ((io_vloadWrites_7_valid && io_flowScalarWrite_valid) && (io_vloadWrites_7_payload_addr == io_flowScalarWrite_payload_addr));
  assign when_WritebackController_l89_334 = ((io_vloadWrites_7_valid && io_flowVectorWrites_0_valid) && (io_vloadWrites_7_payload_addr == io_flowVectorWrites_0_payload_addr));
  assign when_WritebackController_l89_335 = ((io_vloadWrites_7_valid && io_flowVectorWrites_1_valid) && (io_vloadWrites_7_payload_addr == io_flowVectorWrites_1_payload_addr));
  assign when_WritebackController_l89_336 = ((io_vloadWrites_7_valid && io_flowVectorWrites_2_valid) && (io_vloadWrites_7_payload_addr == io_flowVectorWrites_2_payload_addr));
  assign when_WritebackController_l89_337 = ((io_vloadWrites_7_valid && io_flowVectorWrites_3_valid) && (io_vloadWrites_7_payload_addr == io_flowVectorWrites_3_payload_addr));
  assign when_WritebackController_l89_338 = ((io_vloadWrites_7_valid && io_flowVectorWrites_4_valid) && (io_vloadWrites_7_payload_addr == io_flowVectorWrites_4_payload_addr));
  assign when_WritebackController_l89_339 = ((io_vloadWrites_7_valid && io_flowVectorWrites_5_valid) && (io_vloadWrites_7_payload_addr == io_flowVectorWrites_5_payload_addr));
  assign when_WritebackController_l89_340 = ((io_vloadWrites_7_valid && io_flowVectorWrites_6_valid) && (io_vloadWrites_7_payload_addr == io_flowVectorWrites_6_payload_addr));
  assign when_WritebackController_l89_341 = ((io_vloadWrites_7_valid && io_flowVectorWrites_7_valid) && (io_vloadWrites_7_payload_addr == io_flowVectorWrites_7_payload_addr));
  assign when_WritebackController_l89_342 = ((io_flowScalarWrite_valid && io_flowVectorWrites_0_valid) && (io_flowScalarWrite_payload_addr == io_flowVectorWrites_0_payload_addr));
  assign when_WritebackController_l89_343 = ((io_flowScalarWrite_valid && io_flowVectorWrites_1_valid) && (io_flowScalarWrite_payload_addr == io_flowVectorWrites_1_payload_addr));
  assign when_WritebackController_l89_344 = ((io_flowScalarWrite_valid && io_flowVectorWrites_2_valid) && (io_flowScalarWrite_payload_addr == io_flowVectorWrites_2_payload_addr));
  assign when_WritebackController_l89_345 = ((io_flowScalarWrite_valid && io_flowVectorWrites_3_valid) && (io_flowScalarWrite_payload_addr == io_flowVectorWrites_3_payload_addr));
  assign when_WritebackController_l89_346 = ((io_flowScalarWrite_valid && io_flowVectorWrites_4_valid) && (io_flowScalarWrite_payload_addr == io_flowVectorWrites_4_payload_addr));
  assign when_WritebackController_l89_347 = ((io_flowScalarWrite_valid && io_flowVectorWrites_5_valid) && (io_flowScalarWrite_payload_addr == io_flowVectorWrites_5_payload_addr));
  assign when_WritebackController_l89_348 = ((io_flowScalarWrite_valid && io_flowVectorWrites_6_valid) && (io_flowScalarWrite_payload_addr == io_flowVectorWrites_6_payload_addr));
  assign when_WritebackController_l89_349 = ((io_flowScalarWrite_valid && io_flowVectorWrites_7_valid) && (io_flowScalarWrite_payload_addr == io_flowVectorWrites_7_payload_addr));
  assign when_WritebackController_l89_350 = ((io_flowVectorWrites_0_valid && io_flowVectorWrites_1_valid) && (io_flowVectorWrites_0_payload_addr == io_flowVectorWrites_1_payload_addr));
  assign when_WritebackController_l89_351 = ((io_flowVectorWrites_0_valid && io_flowVectorWrites_2_valid) && (io_flowVectorWrites_0_payload_addr == io_flowVectorWrites_2_payload_addr));
  assign when_WritebackController_l89_352 = ((io_flowVectorWrites_0_valid && io_flowVectorWrites_3_valid) && (io_flowVectorWrites_0_payload_addr == io_flowVectorWrites_3_payload_addr));
  assign when_WritebackController_l89_353 = ((io_flowVectorWrites_0_valid && io_flowVectorWrites_4_valid) && (io_flowVectorWrites_0_payload_addr == io_flowVectorWrites_4_payload_addr));
  assign when_WritebackController_l89_354 = ((io_flowVectorWrites_0_valid && io_flowVectorWrites_5_valid) && (io_flowVectorWrites_0_payload_addr == io_flowVectorWrites_5_payload_addr));
  assign when_WritebackController_l89_355 = ((io_flowVectorWrites_0_valid && io_flowVectorWrites_6_valid) && (io_flowVectorWrites_0_payload_addr == io_flowVectorWrites_6_payload_addr));
  assign when_WritebackController_l89_356 = ((io_flowVectorWrites_0_valid && io_flowVectorWrites_7_valid) && (io_flowVectorWrites_0_payload_addr == io_flowVectorWrites_7_payload_addr));
  assign when_WritebackController_l89_357 = ((io_flowVectorWrites_1_valid && io_flowVectorWrites_2_valid) && (io_flowVectorWrites_1_payload_addr == io_flowVectorWrites_2_payload_addr));
  assign when_WritebackController_l89_358 = ((io_flowVectorWrites_1_valid && io_flowVectorWrites_3_valid) && (io_flowVectorWrites_1_payload_addr == io_flowVectorWrites_3_payload_addr));
  assign when_WritebackController_l89_359 = ((io_flowVectorWrites_1_valid && io_flowVectorWrites_4_valid) && (io_flowVectorWrites_1_payload_addr == io_flowVectorWrites_4_payload_addr));
  assign when_WritebackController_l89_360 = ((io_flowVectorWrites_1_valid && io_flowVectorWrites_5_valid) && (io_flowVectorWrites_1_payload_addr == io_flowVectorWrites_5_payload_addr));
  assign when_WritebackController_l89_361 = ((io_flowVectorWrites_1_valid && io_flowVectorWrites_6_valid) && (io_flowVectorWrites_1_payload_addr == io_flowVectorWrites_6_payload_addr));
  assign when_WritebackController_l89_362 = ((io_flowVectorWrites_1_valid && io_flowVectorWrites_7_valid) && (io_flowVectorWrites_1_payload_addr == io_flowVectorWrites_7_payload_addr));
  assign when_WritebackController_l89_363 = ((io_flowVectorWrites_2_valid && io_flowVectorWrites_3_valid) && (io_flowVectorWrites_2_payload_addr == io_flowVectorWrites_3_payload_addr));
  assign when_WritebackController_l89_364 = ((io_flowVectorWrites_2_valid && io_flowVectorWrites_4_valid) && (io_flowVectorWrites_2_payload_addr == io_flowVectorWrites_4_payload_addr));
  assign when_WritebackController_l89_365 = ((io_flowVectorWrites_2_valid && io_flowVectorWrites_5_valid) && (io_flowVectorWrites_2_payload_addr == io_flowVectorWrites_5_payload_addr));
  assign when_WritebackController_l89_366 = ((io_flowVectorWrites_2_valid && io_flowVectorWrites_6_valid) && (io_flowVectorWrites_2_payload_addr == io_flowVectorWrites_6_payload_addr));
  assign when_WritebackController_l89_367 = ((io_flowVectorWrites_2_valid && io_flowVectorWrites_7_valid) && (io_flowVectorWrites_2_payload_addr == io_flowVectorWrites_7_payload_addr));
  assign when_WritebackController_l89_368 = ((io_flowVectorWrites_3_valid && io_flowVectorWrites_4_valid) && (io_flowVectorWrites_3_payload_addr == io_flowVectorWrites_4_payload_addr));
  assign when_WritebackController_l89_369 = ((io_flowVectorWrites_3_valid && io_flowVectorWrites_5_valid) && (io_flowVectorWrites_3_payload_addr == io_flowVectorWrites_5_payload_addr));
  assign when_WritebackController_l89_370 = ((io_flowVectorWrites_3_valid && io_flowVectorWrites_6_valid) && (io_flowVectorWrites_3_payload_addr == io_flowVectorWrites_6_payload_addr));
  assign when_WritebackController_l89_371 = ((io_flowVectorWrites_3_valid && io_flowVectorWrites_7_valid) && (io_flowVectorWrites_3_payload_addr == io_flowVectorWrites_7_payload_addr));
  assign when_WritebackController_l89_372 = ((io_flowVectorWrites_4_valid && io_flowVectorWrites_5_valid) && (io_flowVectorWrites_4_payload_addr == io_flowVectorWrites_5_payload_addr));
  assign when_WritebackController_l89_373 = ((io_flowVectorWrites_4_valid && io_flowVectorWrites_6_valid) && (io_flowVectorWrites_4_payload_addr == io_flowVectorWrites_6_payload_addr));
  assign when_WritebackController_l89_374 = ((io_flowVectorWrites_4_valid && io_flowVectorWrites_7_valid) && (io_flowVectorWrites_4_payload_addr == io_flowVectorWrites_7_payload_addr));
  assign when_WritebackController_l89_375 = ((io_flowVectorWrites_5_valid && io_flowVectorWrites_6_valid) && (io_flowVectorWrites_5_payload_addr == io_flowVectorWrites_6_payload_addr));
  assign when_WritebackController_l89_376 = ((io_flowVectorWrites_5_valid && io_flowVectorWrites_7_valid) && (io_flowVectorWrites_5_payload_addr == io_flowVectorWrites_7_payload_addr));
  assign when_WritebackController_l89_377 = ((io_flowVectorWrites_6_valid && io_flowVectorWrites_7_valid) && (io_flowVectorWrites_6_payload_addr == io_flowVectorWrites_7_payload_addr));
  always @(posedge clk) begin
    if(reset) begin
    end else begin
      if(when_WritebackController_l89) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 0 and port 1 both writing to addr %x", io_aluWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_1) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 0 and port 2 both writing to addr %x", io_aluWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_2) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 0 and port 3 both writing to addr %x", io_aluWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_3) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 0 and port 4 both writing to addr %x", io_aluWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_4) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 0 and port 5 both writing to addr %x", io_aluWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_5) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 0 and port 6 both writing to addr %x", io_aluWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_6) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 0 and port 7 both writing to addr %x", io_aluWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_7) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 0 and port 8 both writing to addr %x", io_aluWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_8) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 0 and port 9 both writing to addr %x", io_aluWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_9) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 0 and port 10 both writing to addr %x", io_aluWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_10) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 0 and port 11 both writing to addr %x", io_aluWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_11) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 0 and port 12 both writing to addr %x", io_aluWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_12) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 0 and port 13 both writing to addr %x", io_aluWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_13) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 0 and port 14 both writing to addr %x", io_aluWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_14) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 0 and port 15 both writing to addr %x", io_aluWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_15) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 0 and port 16 both writing to addr %x", io_aluWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_16) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 0 and port 17 both writing to addr %x", io_aluWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_17) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 0 and port 18 both writing to addr %x", io_aluWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_18) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 0 and port 19 both writing to addr %x", io_aluWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_19) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 0 and port 20 both writing to addr %x", io_aluWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_20) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 0 and port 21 both writing to addr %x", io_aluWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_21) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 0 and port 22 both writing to addr %x", io_aluWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_22) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 0 and port 23 both writing to addr %x", io_aluWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_23) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 0 and port 24 both writing to addr %x", io_aluWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_24) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 0 and port 25 both writing to addr %x", io_aluWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_25) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 0 and port 26 both writing to addr %x", io_aluWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_26) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 0 and port 27 both writing to addr %x", io_aluWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_27) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 1 and port 2 both writing to addr %x", io_valuWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_28) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 1 and port 3 both writing to addr %x", io_valuWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_29) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 1 and port 4 both writing to addr %x", io_valuWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_30) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 1 and port 5 both writing to addr %x", io_valuWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_31) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 1 and port 6 both writing to addr %x", io_valuWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_32) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 1 and port 7 both writing to addr %x", io_valuWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_33) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 1 and port 8 both writing to addr %x", io_valuWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_34) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 1 and port 9 both writing to addr %x", io_valuWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_35) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 1 and port 10 both writing to addr %x", io_valuWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_36) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 1 and port 11 both writing to addr %x", io_valuWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_37) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 1 and port 12 both writing to addr %x", io_valuWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_38) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 1 and port 13 both writing to addr %x", io_valuWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_39) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 1 and port 14 both writing to addr %x", io_valuWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_40) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 1 and port 15 both writing to addr %x", io_valuWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_41) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 1 and port 16 both writing to addr %x", io_valuWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_42) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 1 and port 17 both writing to addr %x", io_valuWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_43) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 1 and port 18 both writing to addr %x", io_valuWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_44) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 1 and port 19 both writing to addr %x", io_valuWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_45) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 1 and port 20 both writing to addr %x", io_valuWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_46) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 1 and port 21 both writing to addr %x", io_valuWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_47) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 1 and port 22 both writing to addr %x", io_valuWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_48) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 1 and port 23 both writing to addr %x", io_valuWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_49) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 1 and port 24 both writing to addr %x", io_valuWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_50) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 1 and port 25 both writing to addr %x", io_valuWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_51) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 1 and port 26 both writing to addr %x", io_valuWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_52) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 1 and port 27 both writing to addr %x", io_valuWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_53) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 2 and port 3 both writing to addr %x", io_valuWrites_1_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_54) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 2 and port 4 both writing to addr %x", io_valuWrites_1_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_55) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 2 and port 5 both writing to addr %x", io_valuWrites_1_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_56) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 2 and port 6 both writing to addr %x", io_valuWrites_1_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_57) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 2 and port 7 both writing to addr %x", io_valuWrites_1_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_58) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 2 and port 8 both writing to addr %x", io_valuWrites_1_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_59) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 2 and port 9 both writing to addr %x", io_valuWrites_1_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_60) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 2 and port 10 both writing to addr %x", io_valuWrites_1_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_61) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 2 and port 11 both writing to addr %x", io_valuWrites_1_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_62) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 2 and port 12 both writing to addr %x", io_valuWrites_1_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_63) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 2 and port 13 both writing to addr %x", io_valuWrites_1_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_64) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 2 and port 14 both writing to addr %x", io_valuWrites_1_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_65) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 2 and port 15 both writing to addr %x", io_valuWrites_1_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_66) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 2 and port 16 both writing to addr %x", io_valuWrites_1_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_67) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 2 and port 17 both writing to addr %x", io_valuWrites_1_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_68) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 2 and port 18 both writing to addr %x", io_valuWrites_1_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_69) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 2 and port 19 both writing to addr %x", io_valuWrites_1_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_70) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 2 and port 20 both writing to addr %x", io_valuWrites_1_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_71) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 2 and port 21 both writing to addr %x", io_valuWrites_1_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_72) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 2 and port 22 both writing to addr %x", io_valuWrites_1_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_73) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 2 and port 23 both writing to addr %x", io_valuWrites_1_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_74) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 2 and port 24 both writing to addr %x", io_valuWrites_1_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_75) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 2 and port 25 both writing to addr %x", io_valuWrites_1_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_76) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 2 and port 26 both writing to addr %x", io_valuWrites_1_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_77) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 2 and port 27 both writing to addr %x", io_valuWrites_1_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_78) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 3 and port 4 both writing to addr %x", io_valuWrites_2_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_79) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 3 and port 5 both writing to addr %x", io_valuWrites_2_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_80) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 3 and port 6 both writing to addr %x", io_valuWrites_2_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_81) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 3 and port 7 both writing to addr %x", io_valuWrites_2_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_82) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 3 and port 8 both writing to addr %x", io_valuWrites_2_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_83) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 3 and port 9 both writing to addr %x", io_valuWrites_2_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_84) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 3 and port 10 both writing to addr %x", io_valuWrites_2_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_85) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 3 and port 11 both writing to addr %x", io_valuWrites_2_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_86) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 3 and port 12 both writing to addr %x", io_valuWrites_2_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_87) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 3 and port 13 both writing to addr %x", io_valuWrites_2_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_88) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 3 and port 14 both writing to addr %x", io_valuWrites_2_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_89) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 3 and port 15 both writing to addr %x", io_valuWrites_2_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_90) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 3 and port 16 both writing to addr %x", io_valuWrites_2_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_91) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 3 and port 17 both writing to addr %x", io_valuWrites_2_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_92) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 3 and port 18 both writing to addr %x", io_valuWrites_2_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_93) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 3 and port 19 both writing to addr %x", io_valuWrites_2_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_94) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 3 and port 20 both writing to addr %x", io_valuWrites_2_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_95) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 3 and port 21 both writing to addr %x", io_valuWrites_2_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_96) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 3 and port 22 both writing to addr %x", io_valuWrites_2_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_97) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 3 and port 23 both writing to addr %x", io_valuWrites_2_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_98) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 3 and port 24 both writing to addr %x", io_valuWrites_2_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_99) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 3 and port 25 both writing to addr %x", io_valuWrites_2_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_100) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 3 and port 26 both writing to addr %x", io_valuWrites_2_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_101) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 3 and port 27 both writing to addr %x", io_valuWrites_2_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_102) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 4 and port 5 both writing to addr %x", io_valuWrites_3_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_103) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 4 and port 6 both writing to addr %x", io_valuWrites_3_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_104) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 4 and port 7 both writing to addr %x", io_valuWrites_3_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_105) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 4 and port 8 both writing to addr %x", io_valuWrites_3_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_106) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 4 and port 9 both writing to addr %x", io_valuWrites_3_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_107) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 4 and port 10 both writing to addr %x", io_valuWrites_3_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_108) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 4 and port 11 both writing to addr %x", io_valuWrites_3_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_109) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 4 and port 12 both writing to addr %x", io_valuWrites_3_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_110) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 4 and port 13 both writing to addr %x", io_valuWrites_3_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_111) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 4 and port 14 both writing to addr %x", io_valuWrites_3_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_112) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 4 and port 15 both writing to addr %x", io_valuWrites_3_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_113) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 4 and port 16 both writing to addr %x", io_valuWrites_3_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_114) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 4 and port 17 both writing to addr %x", io_valuWrites_3_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_115) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 4 and port 18 both writing to addr %x", io_valuWrites_3_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_116) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 4 and port 19 both writing to addr %x", io_valuWrites_3_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_117) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 4 and port 20 both writing to addr %x", io_valuWrites_3_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_118) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 4 and port 21 both writing to addr %x", io_valuWrites_3_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_119) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 4 and port 22 both writing to addr %x", io_valuWrites_3_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_120) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 4 and port 23 both writing to addr %x", io_valuWrites_3_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_121) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 4 and port 24 both writing to addr %x", io_valuWrites_3_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_122) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 4 and port 25 both writing to addr %x", io_valuWrites_3_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_123) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 4 and port 26 both writing to addr %x", io_valuWrites_3_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_124) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 4 and port 27 both writing to addr %x", io_valuWrites_3_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_125) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 5 and port 6 both writing to addr %x", io_valuWrites_4_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_126) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 5 and port 7 both writing to addr %x", io_valuWrites_4_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_127) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 5 and port 8 both writing to addr %x", io_valuWrites_4_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_128) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 5 and port 9 both writing to addr %x", io_valuWrites_4_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_129) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 5 and port 10 both writing to addr %x", io_valuWrites_4_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_130) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 5 and port 11 both writing to addr %x", io_valuWrites_4_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_131) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 5 and port 12 both writing to addr %x", io_valuWrites_4_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_132) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 5 and port 13 both writing to addr %x", io_valuWrites_4_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_133) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 5 and port 14 both writing to addr %x", io_valuWrites_4_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_134) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 5 and port 15 both writing to addr %x", io_valuWrites_4_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_135) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 5 and port 16 both writing to addr %x", io_valuWrites_4_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_136) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 5 and port 17 both writing to addr %x", io_valuWrites_4_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_137) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 5 and port 18 both writing to addr %x", io_valuWrites_4_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_138) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 5 and port 19 both writing to addr %x", io_valuWrites_4_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_139) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 5 and port 20 both writing to addr %x", io_valuWrites_4_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_140) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 5 and port 21 both writing to addr %x", io_valuWrites_4_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_141) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 5 and port 22 both writing to addr %x", io_valuWrites_4_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_142) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 5 and port 23 both writing to addr %x", io_valuWrites_4_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_143) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 5 and port 24 both writing to addr %x", io_valuWrites_4_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_144) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 5 and port 25 both writing to addr %x", io_valuWrites_4_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_145) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 5 and port 26 both writing to addr %x", io_valuWrites_4_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_146) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 5 and port 27 both writing to addr %x", io_valuWrites_4_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_147) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 6 and port 7 both writing to addr %x", io_valuWrites_5_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_148) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 6 and port 8 both writing to addr %x", io_valuWrites_5_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_149) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 6 and port 9 both writing to addr %x", io_valuWrites_5_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_150) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 6 and port 10 both writing to addr %x", io_valuWrites_5_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_151) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 6 and port 11 both writing to addr %x", io_valuWrites_5_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_152) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 6 and port 12 both writing to addr %x", io_valuWrites_5_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_153) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 6 and port 13 both writing to addr %x", io_valuWrites_5_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_154) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 6 and port 14 both writing to addr %x", io_valuWrites_5_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_155) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 6 and port 15 both writing to addr %x", io_valuWrites_5_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_156) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 6 and port 16 both writing to addr %x", io_valuWrites_5_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_157) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 6 and port 17 both writing to addr %x", io_valuWrites_5_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_158) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 6 and port 18 both writing to addr %x", io_valuWrites_5_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_159) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 6 and port 19 both writing to addr %x", io_valuWrites_5_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_160) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 6 and port 20 both writing to addr %x", io_valuWrites_5_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_161) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 6 and port 21 both writing to addr %x", io_valuWrites_5_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_162) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 6 and port 22 both writing to addr %x", io_valuWrites_5_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_163) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 6 and port 23 both writing to addr %x", io_valuWrites_5_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_164) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 6 and port 24 both writing to addr %x", io_valuWrites_5_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_165) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 6 and port 25 both writing to addr %x", io_valuWrites_5_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_166) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 6 and port 26 both writing to addr %x", io_valuWrites_5_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_167) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 6 and port 27 both writing to addr %x", io_valuWrites_5_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_168) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 7 and port 8 both writing to addr %x", io_valuWrites_6_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_169) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 7 and port 9 both writing to addr %x", io_valuWrites_6_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_170) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 7 and port 10 both writing to addr %x", io_valuWrites_6_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_171) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 7 and port 11 both writing to addr %x", io_valuWrites_6_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_172) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 7 and port 12 both writing to addr %x", io_valuWrites_6_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_173) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 7 and port 13 both writing to addr %x", io_valuWrites_6_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_174) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 7 and port 14 both writing to addr %x", io_valuWrites_6_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_175) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 7 and port 15 both writing to addr %x", io_valuWrites_6_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_176) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 7 and port 16 both writing to addr %x", io_valuWrites_6_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_177) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 7 and port 17 both writing to addr %x", io_valuWrites_6_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_178) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 7 and port 18 both writing to addr %x", io_valuWrites_6_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_179) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 7 and port 19 both writing to addr %x", io_valuWrites_6_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_180) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 7 and port 20 both writing to addr %x", io_valuWrites_6_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_181) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 7 and port 21 both writing to addr %x", io_valuWrites_6_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_182) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 7 and port 22 both writing to addr %x", io_valuWrites_6_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_183) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 7 and port 23 both writing to addr %x", io_valuWrites_6_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_184) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 7 and port 24 both writing to addr %x", io_valuWrites_6_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_185) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 7 and port 25 both writing to addr %x", io_valuWrites_6_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_186) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 7 and port 26 both writing to addr %x", io_valuWrites_6_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_187) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 7 and port 27 both writing to addr %x", io_valuWrites_6_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_188) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 8 and port 9 both writing to addr %x", io_valuWrites_7_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_189) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 8 and port 10 both writing to addr %x", io_valuWrites_7_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_190) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 8 and port 11 both writing to addr %x", io_valuWrites_7_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_191) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 8 and port 12 both writing to addr %x", io_valuWrites_7_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_192) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 8 and port 13 both writing to addr %x", io_valuWrites_7_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_193) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 8 and port 14 both writing to addr %x", io_valuWrites_7_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_194) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 8 and port 15 both writing to addr %x", io_valuWrites_7_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_195) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 8 and port 16 both writing to addr %x", io_valuWrites_7_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_196) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 8 and port 17 both writing to addr %x", io_valuWrites_7_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_197) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 8 and port 18 both writing to addr %x", io_valuWrites_7_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_198) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 8 and port 19 both writing to addr %x", io_valuWrites_7_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_199) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 8 and port 20 both writing to addr %x", io_valuWrites_7_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_200) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 8 and port 21 both writing to addr %x", io_valuWrites_7_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_201) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 8 and port 22 both writing to addr %x", io_valuWrites_7_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_202) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 8 and port 23 both writing to addr %x", io_valuWrites_7_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_203) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 8 and port 24 both writing to addr %x", io_valuWrites_7_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_204) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 8 and port 25 both writing to addr %x", io_valuWrites_7_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_205) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 8 and port 26 both writing to addr %x", io_valuWrites_7_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_206) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 8 and port 27 both writing to addr %x", io_valuWrites_7_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_207) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 9 and port 10 both writing to addr %x", io_loadWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_208) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 9 and port 11 both writing to addr %x", io_loadWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_209) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 9 and port 12 both writing to addr %x", io_loadWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_210) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 9 and port 13 both writing to addr %x", io_loadWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_211) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 9 and port 14 both writing to addr %x", io_loadWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_212) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 9 and port 15 both writing to addr %x", io_loadWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_213) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 9 and port 16 both writing to addr %x", io_loadWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_214) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 9 and port 17 both writing to addr %x", io_loadWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_215) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 9 and port 18 both writing to addr %x", io_loadWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_216) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 9 and port 19 both writing to addr %x", io_loadWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_217) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 9 and port 20 both writing to addr %x", io_loadWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_218) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 9 and port 21 both writing to addr %x", io_loadWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_219) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 9 and port 22 both writing to addr %x", io_loadWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_220) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 9 and port 23 both writing to addr %x", io_loadWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_221) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 9 and port 24 both writing to addr %x", io_loadWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_222) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 9 and port 25 both writing to addr %x", io_loadWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_223) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 9 and port 26 both writing to addr %x", io_loadWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_224) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 9 and port 27 both writing to addr %x", io_loadWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_225) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 10 and port 11 both writing to addr %x", io_constWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_226) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 10 and port 12 both writing to addr %x", io_constWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_227) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 10 and port 13 both writing to addr %x", io_constWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_228) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 10 and port 14 both writing to addr %x", io_constWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_229) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 10 and port 15 both writing to addr %x", io_constWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_230) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 10 and port 16 both writing to addr %x", io_constWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_231) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 10 and port 17 both writing to addr %x", io_constWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_232) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 10 and port 18 both writing to addr %x", io_constWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_233) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 10 and port 19 both writing to addr %x", io_constWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_234) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 10 and port 20 both writing to addr %x", io_constWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_235) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 10 and port 21 both writing to addr %x", io_constWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_236) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 10 and port 22 both writing to addr %x", io_constWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_237) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 10 and port 23 both writing to addr %x", io_constWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_238) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 10 and port 24 both writing to addr %x", io_constWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_239) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 10 and port 25 both writing to addr %x", io_constWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_240) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 10 and port 26 both writing to addr %x", io_constWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_241) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 10 and port 27 both writing to addr %x", io_constWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_242) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 11 and port 12 both writing to addr %x", io_vloadWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_243) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 11 and port 13 both writing to addr %x", io_vloadWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_244) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 11 and port 14 both writing to addr %x", io_vloadWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_245) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 11 and port 15 both writing to addr %x", io_vloadWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_246) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 11 and port 16 both writing to addr %x", io_vloadWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_247) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 11 and port 17 both writing to addr %x", io_vloadWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_248) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 11 and port 18 both writing to addr %x", io_vloadWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_249) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 11 and port 19 both writing to addr %x", io_vloadWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_250) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 11 and port 20 both writing to addr %x", io_vloadWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_251) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 11 and port 21 both writing to addr %x", io_vloadWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_252) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 11 and port 22 both writing to addr %x", io_vloadWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_253) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 11 and port 23 both writing to addr %x", io_vloadWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_254) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 11 and port 24 both writing to addr %x", io_vloadWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_255) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 11 and port 25 both writing to addr %x", io_vloadWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_256) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 11 and port 26 both writing to addr %x", io_vloadWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_257) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 11 and port 27 both writing to addr %x", io_vloadWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_258) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 12 and port 13 both writing to addr %x", io_vloadWrites_1_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_259) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 12 and port 14 both writing to addr %x", io_vloadWrites_1_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_260) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 12 and port 15 both writing to addr %x", io_vloadWrites_1_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_261) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 12 and port 16 both writing to addr %x", io_vloadWrites_1_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_262) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 12 and port 17 both writing to addr %x", io_vloadWrites_1_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_263) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 12 and port 18 both writing to addr %x", io_vloadWrites_1_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_264) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 12 and port 19 both writing to addr %x", io_vloadWrites_1_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_265) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 12 and port 20 both writing to addr %x", io_vloadWrites_1_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_266) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 12 and port 21 both writing to addr %x", io_vloadWrites_1_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_267) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 12 and port 22 both writing to addr %x", io_vloadWrites_1_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_268) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 12 and port 23 both writing to addr %x", io_vloadWrites_1_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_269) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 12 and port 24 both writing to addr %x", io_vloadWrites_1_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_270) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 12 and port 25 both writing to addr %x", io_vloadWrites_1_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_271) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 12 and port 26 both writing to addr %x", io_vloadWrites_1_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_272) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 12 and port 27 both writing to addr %x", io_vloadWrites_1_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_273) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 13 and port 14 both writing to addr %x", io_vloadWrites_2_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_274) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 13 and port 15 both writing to addr %x", io_vloadWrites_2_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_275) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 13 and port 16 both writing to addr %x", io_vloadWrites_2_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_276) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 13 and port 17 both writing to addr %x", io_vloadWrites_2_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_277) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 13 and port 18 both writing to addr %x", io_vloadWrites_2_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_278) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 13 and port 19 both writing to addr %x", io_vloadWrites_2_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_279) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 13 and port 20 both writing to addr %x", io_vloadWrites_2_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_280) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 13 and port 21 both writing to addr %x", io_vloadWrites_2_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_281) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 13 and port 22 both writing to addr %x", io_vloadWrites_2_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_282) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 13 and port 23 both writing to addr %x", io_vloadWrites_2_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_283) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 13 and port 24 both writing to addr %x", io_vloadWrites_2_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_284) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 13 and port 25 both writing to addr %x", io_vloadWrites_2_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_285) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 13 and port 26 both writing to addr %x", io_vloadWrites_2_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_286) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 13 and port 27 both writing to addr %x", io_vloadWrites_2_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_287) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 14 and port 15 both writing to addr %x", io_vloadWrites_3_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_288) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 14 and port 16 both writing to addr %x", io_vloadWrites_3_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_289) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 14 and port 17 both writing to addr %x", io_vloadWrites_3_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_290) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 14 and port 18 both writing to addr %x", io_vloadWrites_3_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_291) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 14 and port 19 both writing to addr %x", io_vloadWrites_3_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_292) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 14 and port 20 both writing to addr %x", io_vloadWrites_3_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_293) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 14 and port 21 both writing to addr %x", io_vloadWrites_3_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_294) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 14 and port 22 both writing to addr %x", io_vloadWrites_3_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_295) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 14 and port 23 both writing to addr %x", io_vloadWrites_3_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_296) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 14 and port 24 both writing to addr %x", io_vloadWrites_3_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_297) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 14 and port 25 both writing to addr %x", io_vloadWrites_3_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_298) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 14 and port 26 both writing to addr %x", io_vloadWrites_3_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_299) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 14 and port 27 both writing to addr %x", io_vloadWrites_3_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_300) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 15 and port 16 both writing to addr %x", io_vloadWrites_4_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_301) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 15 and port 17 both writing to addr %x", io_vloadWrites_4_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_302) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 15 and port 18 both writing to addr %x", io_vloadWrites_4_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_303) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 15 and port 19 both writing to addr %x", io_vloadWrites_4_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_304) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 15 and port 20 both writing to addr %x", io_vloadWrites_4_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_305) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 15 and port 21 both writing to addr %x", io_vloadWrites_4_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_306) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 15 and port 22 both writing to addr %x", io_vloadWrites_4_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_307) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 15 and port 23 both writing to addr %x", io_vloadWrites_4_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_308) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 15 and port 24 both writing to addr %x", io_vloadWrites_4_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_309) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 15 and port 25 both writing to addr %x", io_vloadWrites_4_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_310) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 15 and port 26 both writing to addr %x", io_vloadWrites_4_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_311) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 15 and port 27 both writing to addr %x", io_vloadWrites_4_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_312) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 16 and port 17 both writing to addr %x", io_vloadWrites_5_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_313) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 16 and port 18 both writing to addr %x", io_vloadWrites_5_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_314) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 16 and port 19 both writing to addr %x", io_vloadWrites_5_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_315) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 16 and port 20 both writing to addr %x", io_vloadWrites_5_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_316) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 16 and port 21 both writing to addr %x", io_vloadWrites_5_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_317) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 16 and port 22 both writing to addr %x", io_vloadWrites_5_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_318) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 16 and port 23 both writing to addr %x", io_vloadWrites_5_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_319) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 16 and port 24 both writing to addr %x", io_vloadWrites_5_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_320) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 16 and port 25 both writing to addr %x", io_vloadWrites_5_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_321) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 16 and port 26 both writing to addr %x", io_vloadWrites_5_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_322) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 16 and port 27 both writing to addr %x", io_vloadWrites_5_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_323) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 17 and port 18 both writing to addr %x", io_vloadWrites_6_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_324) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 17 and port 19 both writing to addr %x", io_vloadWrites_6_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_325) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 17 and port 20 both writing to addr %x", io_vloadWrites_6_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_326) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 17 and port 21 both writing to addr %x", io_vloadWrites_6_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_327) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 17 and port 22 both writing to addr %x", io_vloadWrites_6_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_328) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 17 and port 23 both writing to addr %x", io_vloadWrites_6_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_329) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 17 and port 24 both writing to addr %x", io_vloadWrites_6_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_330) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 17 and port 25 both writing to addr %x", io_vloadWrites_6_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_331) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 17 and port 26 both writing to addr %x", io_vloadWrites_6_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_332) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 17 and port 27 both writing to addr %x", io_vloadWrites_6_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_333) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 18 and port 19 both writing to addr %x", io_vloadWrites_7_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_334) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 18 and port 20 both writing to addr %x", io_vloadWrites_7_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_335) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 18 and port 21 both writing to addr %x", io_vloadWrites_7_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_336) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 18 and port 22 both writing to addr %x", io_vloadWrites_7_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_337) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 18 and port 23 both writing to addr %x", io_vloadWrites_7_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_338) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 18 and port 24 both writing to addr %x", io_vloadWrites_7_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_339) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 18 and port 25 both writing to addr %x", io_vloadWrites_7_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_340) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 18 and port 26 both writing to addr %x", io_vloadWrites_7_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_341) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 18 and port 27 both writing to addr %x", io_vloadWrites_7_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_342) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 19 and port 20 both writing to addr %x", io_flowScalarWrite_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_343) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 19 and port 21 both writing to addr %x", io_flowScalarWrite_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_344) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 19 and port 22 both writing to addr %x", io_flowScalarWrite_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_345) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 19 and port 23 both writing to addr %x", io_flowScalarWrite_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_346) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 19 and port 24 both writing to addr %x", io_flowScalarWrite_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_347) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 19 and port 25 both writing to addr %x", io_flowScalarWrite_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_348) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 19 and port 26 both writing to addr %x", io_flowScalarWrite_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_349) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 19 and port 27 both writing to addr %x", io_flowScalarWrite_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_350) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 20 and port 21 both writing to addr %x", io_flowVectorWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_351) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 20 and port 22 both writing to addr %x", io_flowVectorWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_352) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 20 and port 23 both writing to addr %x", io_flowVectorWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_353) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 20 and port 24 both writing to addr %x", io_flowVectorWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_354) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 20 and port 25 both writing to addr %x", io_flowVectorWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_355) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 20 and port 26 both writing to addr %x", io_flowVectorWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_356) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 20 and port 27 both writing to addr %x", io_flowVectorWrites_0_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_357) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 21 and port 22 both writing to addr %x", io_flowVectorWrites_1_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_358) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 21 and port 23 both writing to addr %x", io_flowVectorWrites_1_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_359) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 21 and port 24 both writing to addr %x", io_flowVectorWrites_1_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_360) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 21 and port 25 both writing to addr %x", io_flowVectorWrites_1_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_361) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 21 and port 26 both writing to addr %x", io_flowVectorWrites_1_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_362) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 21 and port 27 both writing to addr %x", io_flowVectorWrites_1_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_363) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 22 and port 23 both writing to addr %x", io_flowVectorWrites_2_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_364) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 22 and port 24 both writing to addr %x", io_flowVectorWrites_2_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_365) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 22 and port 25 both writing to addr %x", io_flowVectorWrites_2_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_366) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 22 and port 26 both writing to addr %x", io_flowVectorWrites_2_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_367) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 22 and port 27 both writing to addr %x", io_flowVectorWrites_2_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_368) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 23 and port 24 both writing to addr %x", io_flowVectorWrites_3_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_369) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 23 and port 25 both writing to addr %x", io_flowVectorWrites_3_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_370) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 23 and port 26 both writing to addr %x", io_flowVectorWrites_3_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_371) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 23 and port 27 both writing to addr %x", io_flowVectorWrites_3_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_372) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 24 and port 25 both writing to addr %x", io_flowVectorWrites_4_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_373) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 24 and port 26 both writing to addr %x", io_flowVectorWrites_4_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_374) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 24 and port 27 both writing to addr %x", io_flowVectorWrites_4_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_375) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 25 and port 26 both writing to addr %x", io_flowVectorWrites_5_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_376) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 25 and port 27 both writing to addr %x", io_flowVectorWrites_5_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
      if(when_WritebackController_l89_377) begin
        `ifndef SYNTHESIS
          `ifdef FORMAL
            assert(1'b0); // core.scala:L522
          `else
            if(!1'b0) begin
              $display("NOTE WAW CONFLICT detected: port 26 and port 27 both writing to addr %x", io_flowVectorWrites_6_payload_addr); // core.scala:L522
            end
          `endif
        `endif
      end
    end
  end


endmodule
