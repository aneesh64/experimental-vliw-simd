// Generator : SpinalHDL v1.10.2a    git head : a348a60b7e8b6a455c72e1536ec3d74a2ea16935
// Component : MemoryEngine
// Git hash  : 2b1c34e10fcfebdb7017c9a507f6d279f35a00fa

`timescale 1ns/1ps

module MemoryEngine (
  input  wire          io_loadSlots_0_valid,
  input  wire [2:0]    io_loadSlots_0_opcode,
  input  wire [10:0]   io_loadSlots_0_dest,
  input  wire [10:0]   io_loadSlots_0_addrReg,
  input  wire [2:0]    io_loadSlots_0_offset,
  input  wire [31:0]   io_loadSlots_0_immediate,
  input  wire          io_storeSlots_0_valid,
  input  wire [1:0]    io_storeSlots_0_opcode,
  input  wire [10:0]   io_storeSlots_0_addrReg,
  input  wire [10:0]   io_storeSlots_0_srcReg,
  input  wire          io_valid,
  input  wire [31:0]   io_loadAddrData_0,
  input  wire [31:0]   io_storeAddrData_0,
  input  wire [31:0]   io_storeSrcData_0,
  input  wire [31:0]   io_vstoreSrcData_0_0,
  input  wire [31:0]   io_vstoreSrcData_0_1,
  input  wire [31:0]   io_vstoreSrcData_0_2,
  input  wire [31:0]   io_vstoreSrcData_0_3,
  input  wire [31:0]   io_vstoreSrcData_0_4,
  input  wire [31:0]   io_vstoreSrcData_0_5,
  input  wire [31:0]   io_vstoreSrcData_0_6,
  input  wire [31:0]   io_vstoreSrcData_0_7,
  output reg           io_axiMaster_aw_valid,
  input  wire          io_axiMaster_aw_ready,
  output reg  [31:0]   io_axiMaster_aw_payload_addr,
  output wire [3:0]    io_axiMaster_aw_payload_id,
  output reg  [7:0]    io_axiMaster_aw_payload_len,
  output reg  [2:0]    io_axiMaster_aw_payload_size,
  output wire [1:0]    io_axiMaster_aw_payload_burst,
  output reg           io_axiMaster_w_valid,
  input  wire          io_axiMaster_w_ready,
  output reg  [511:0]  io_axiMaster_w_payload_data,
  output reg  [63:0]   io_axiMaster_w_payload_strb,
  output reg           io_axiMaster_w_payload_last,
  input  wire          io_axiMaster_b_valid,
  output reg           io_axiMaster_b_ready,
  input  wire [3:0]    io_axiMaster_b_payload_id,
  input  wire [1:0]    io_axiMaster_b_payload_resp,
  output wire          io_axiMaster_ar_valid,
  input  wire          io_axiMaster_ar_ready,
  output wire [31:0]   io_axiMaster_ar_payload_addr,
  output wire [3:0]    io_axiMaster_ar_payload_id,
  output wire [7:0]    io_axiMaster_ar_payload_len,
  output wire [2:0]    io_axiMaster_ar_payload_size,
  output wire [1:0]    io_axiMaster_ar_payload_burst,
  input  wire          io_axiMaster_r_valid,
  output wire          io_axiMaster_r_ready,
  input  wire [511:0]  io_axiMaster_r_payload_data,
  input  wire [3:0]    io_axiMaster_r_payload_id,
  input  wire [1:0]    io_axiMaster_r_payload_resp,
  input  wire          io_axiMaster_r_payload_last,
  output reg           io_loadWriteReqs_0_valid,
  output reg  [10:0]   io_loadWriteReqs_0_payload_addr,
  output reg  [31:0]   io_loadWriteReqs_0_payload_data,
  output reg           io_constWriteReqs_0_valid,
  output reg  [10:0]   io_constWriteReqs_0_payload_addr,
  output reg  [31:0]   io_constWriteReqs_0_payload_data,
  output reg           io_vloadWriteReqs_0_0_valid,
  output reg  [10:0]   io_vloadWriteReqs_0_0_payload_addr,
  output reg  [31:0]   io_vloadWriteReqs_0_0_payload_data,
  output reg           io_vloadWriteReqs_0_1_valid,
  output reg  [10:0]   io_vloadWriteReqs_0_1_payload_addr,
  output reg  [31:0]   io_vloadWriteReqs_0_1_payload_data,
  output reg           io_vloadWriteReqs_0_2_valid,
  output reg  [10:0]   io_vloadWriteReqs_0_2_payload_addr,
  output reg  [31:0]   io_vloadWriteReqs_0_2_payload_data,
  output reg           io_vloadWriteReqs_0_3_valid,
  output reg  [10:0]   io_vloadWriteReqs_0_3_payload_addr,
  output reg  [31:0]   io_vloadWriteReqs_0_3_payload_data,
  output reg           io_vloadWriteReqs_0_4_valid,
  output reg  [10:0]   io_vloadWriteReqs_0_4_payload_addr,
  output reg  [31:0]   io_vloadWriteReqs_0_4_payload_data,
  output reg           io_vloadWriteReqs_0_5_valid,
  output reg  [10:0]   io_vloadWriteReqs_0_5_payload_addr,
  output reg  [31:0]   io_vloadWriteReqs_0_5_payload_data,
  output reg           io_vloadWriteReqs_0_6_valid,
  output reg  [10:0]   io_vloadWriteReqs_0_6_payload_addr,
  output reg  [31:0]   io_vloadWriteReqs_0_6_payload_data,
  output reg           io_vloadWriteReqs_0_7_valid,
  output reg  [10:0]   io_vloadWriteReqs_0_7_payload_addr,
  output reg  [31:0]   io_vloadWriteReqs_0_7_payload_data,
  output reg           io_stall,
  input  wire          clk,
  input  wire          reset
);
  localparam MemState_IDLE = 2'd0;
  localparam MemState_STORE_AW_W = 2'd1;
  localparam MemState_STORE_B = 2'd2;

  reg                 storeReqFifo_io_push_valid;
  reg        [31:0]   storeReqFifo_io_push_payload_axiAddr;
  reg        [511:0]  storeReqFifo_io_push_payload_wdata;
  reg        [63:0]   storeReqFifo_io_push_payload_wstrb;
  reg                 storeReqFifo_io_pop_ready;
  wire                storeReqFifo_io_push_ready;
  wire                storeReqFifo_io_pop_valid;
  wire       [31:0]   storeReqFifo_io_pop_payload_axiAddr;
  wire       [511:0]  storeReqFifo_io_pop_payload_wdata;
  wire       [63:0]   storeReqFifo_io_pop_payload_wstrb;
  wire       [3:0]    storeReqFifo_io_occupancy;
  wire       [3:0]    storeReqFifo_io_availability;
  wire       [33:0]   _zz__zz_loadReqEntry_wordOff;
  wire       [29:0]   _zz_loadReqEntry_wordOff_1;
  wire       [33:0]   _zz__zz_loadReqEntry_axiAddr_2;
  wire       [31:0]   _zz__zz_loadReqEntry_axiAddr_2_1;
  wire       [31:0]   _zz__zz_loadReqEntry_axiAddr_2_2;
  wire       [10:0]   _zz_loadReqEntry_destAddr;
  wire       [29:0]   _zz_loadReqEntry_wordOff_2;
  wire       [33:0]   _zz__zz_io_push_payload_axiAddr_1;
  wire       [29:0]   _zz__zz_when_MemoryEngine_l235;
  wire       [2:0]    axiSizeVal;
  wire                when_MemoryEngine_l103;
  wire       [607:0]  _zz_io_push_payload_axiAddr;
  reg                 loadReqValid;
  reg        [31:0]   loadReqEntry_axiAddr;
  reg        [10:0]   loadReqEntry_destAddr;
  reg                 loadReqEntry_isVector;
  reg        [0:0]    loadReqEntry_slotIdx;
  reg        [3:0]    loadReqEntry_wordOff;
  reg                 anyLoadOp;
  wire                isLoadOp_0;
  reg                 anyStoreOp;
  wire                isStoreOp_0;
  wire                when_MemoryEngine_l167;
  wire                when_MemoryEngine_l172;
  wire                when_MemoryEngine_l180;
  wire       [31:0]   _zz_loadReqEntry_wordOff;
  wire       [31:0]   _zz_loadReqEntry_axiAddr;
  wire       [31:0]   _zz_loadReqEntry_axiAddr_1;
  wire       [31:0]   _zz_loadReqEntry_axiAddr_2;
  wire                when_MemoryEngine_l215;
  wire       [31:0]   _zz_io_push_payload_axiAddr_1;
  wire       [3:0]    _zz_when_MemoryEngine_l235;
  reg        [511:0]  _zz_io_push_payload_wdata;
  reg        [63:0]   _zz_io_push_payload_wstrb;
  wire                when_MemoryEngine_l235;
  wire                when_MemoryEngine_l235_1;
  wire                when_MemoryEngine_l235_2;
  wire                when_MemoryEngine_l235_3;
  wire                when_MemoryEngine_l235_4;
  wire                when_MemoryEngine_l235_5;
  wire                when_MemoryEngine_l235_6;
  wire                when_MemoryEngine_l235_7;
  wire                when_MemoryEngine_l235_8;
  wire                when_MemoryEngine_l235_9;
  wire                when_MemoryEngine_l235_10;
  wire                when_MemoryEngine_l235_11;
  wire                when_MemoryEngine_l235_12;
  wire                when_MemoryEngine_l235_13;
  wire                when_MemoryEngine_l235_14;
  wire                when_MemoryEngine_l235_15;
  wire       [3:0]    _zz_when_MemoryEngine_l246;
  wire                when_MemoryEngine_l246;
  wire                when_MemoryEngine_l246_1;
  wire                when_MemoryEngine_l246_2;
  wire                when_MemoryEngine_l246_3;
  wire                when_MemoryEngine_l246_4;
  wire                when_MemoryEngine_l246_5;
  wire                when_MemoryEngine_l246_6;
  wire                when_MemoryEngine_l246_7;
  wire                when_MemoryEngine_l246_8;
  wire                when_MemoryEngine_l246_9;
  wire                when_MemoryEngine_l246_10;
  wire                when_MemoryEngine_l246_11;
  wire                when_MemoryEngine_l246_12;
  wire                when_MemoryEngine_l246_13;
  wire                when_MemoryEngine_l246_14;
  wire                when_MemoryEngine_l246_15;
  wire       [3:0]    _zz_when_MemoryEngine_l246_1;
  wire                when_MemoryEngine_l246_16;
  wire                when_MemoryEngine_l246_17;
  wire                when_MemoryEngine_l246_18;
  wire                when_MemoryEngine_l246_19;
  wire                when_MemoryEngine_l246_20;
  wire                when_MemoryEngine_l246_21;
  wire                when_MemoryEngine_l246_22;
  wire                when_MemoryEngine_l246_23;
  wire                when_MemoryEngine_l246_24;
  wire                when_MemoryEngine_l246_25;
  wire                when_MemoryEngine_l246_26;
  wire                when_MemoryEngine_l246_27;
  wire                when_MemoryEngine_l246_28;
  wire                when_MemoryEngine_l246_29;
  wire                when_MemoryEngine_l246_30;
  wire                when_MemoryEngine_l246_31;
  wire       [3:0]    _zz_when_MemoryEngine_l246_2;
  wire                when_MemoryEngine_l246_32;
  wire                when_MemoryEngine_l246_33;
  wire                when_MemoryEngine_l246_34;
  wire                when_MemoryEngine_l246_35;
  wire                when_MemoryEngine_l246_36;
  wire                when_MemoryEngine_l246_37;
  wire                when_MemoryEngine_l246_38;
  wire                when_MemoryEngine_l246_39;
  wire                when_MemoryEngine_l246_40;
  wire                when_MemoryEngine_l246_41;
  wire                when_MemoryEngine_l246_42;
  wire                when_MemoryEngine_l246_43;
  wire                when_MemoryEngine_l246_44;
  wire                when_MemoryEngine_l246_45;
  wire                when_MemoryEngine_l246_46;
  wire                when_MemoryEngine_l246_47;
  wire       [3:0]    _zz_when_MemoryEngine_l246_3;
  wire                when_MemoryEngine_l246_48;
  wire                when_MemoryEngine_l246_49;
  wire                when_MemoryEngine_l246_50;
  wire                when_MemoryEngine_l246_51;
  wire                when_MemoryEngine_l246_52;
  wire                when_MemoryEngine_l246_53;
  wire                when_MemoryEngine_l246_54;
  wire                when_MemoryEngine_l246_55;
  wire                when_MemoryEngine_l246_56;
  wire                when_MemoryEngine_l246_57;
  wire                when_MemoryEngine_l246_58;
  wire                when_MemoryEngine_l246_59;
  wire                when_MemoryEngine_l246_60;
  wire                when_MemoryEngine_l246_61;
  wire                when_MemoryEngine_l246_62;
  wire                when_MemoryEngine_l246_63;
  wire       [3:0]    _zz_when_MemoryEngine_l246_4;
  wire                when_MemoryEngine_l246_64;
  wire                when_MemoryEngine_l246_65;
  wire                when_MemoryEngine_l246_66;
  wire                when_MemoryEngine_l246_67;
  wire                when_MemoryEngine_l246_68;
  wire                when_MemoryEngine_l246_69;
  wire                when_MemoryEngine_l246_70;
  wire                when_MemoryEngine_l246_71;
  wire                when_MemoryEngine_l246_72;
  wire                when_MemoryEngine_l246_73;
  wire                when_MemoryEngine_l246_74;
  wire                when_MemoryEngine_l246_75;
  wire                when_MemoryEngine_l246_76;
  wire                when_MemoryEngine_l246_77;
  wire                when_MemoryEngine_l246_78;
  wire                when_MemoryEngine_l246_79;
  wire       [3:0]    _zz_when_MemoryEngine_l246_5;
  wire                when_MemoryEngine_l246_80;
  wire                when_MemoryEngine_l246_81;
  wire                when_MemoryEngine_l246_82;
  wire                when_MemoryEngine_l246_83;
  wire                when_MemoryEngine_l246_84;
  wire                when_MemoryEngine_l246_85;
  wire                when_MemoryEngine_l246_86;
  wire                when_MemoryEngine_l246_87;
  wire                when_MemoryEngine_l246_88;
  wire                when_MemoryEngine_l246_89;
  wire                when_MemoryEngine_l246_90;
  wire                when_MemoryEngine_l246_91;
  wire                when_MemoryEngine_l246_92;
  wire                when_MemoryEngine_l246_93;
  wire                when_MemoryEngine_l246_94;
  wire                when_MemoryEngine_l246_95;
  wire       [3:0]    _zz_when_MemoryEngine_l246_6;
  wire                when_MemoryEngine_l246_96;
  wire                when_MemoryEngine_l246_97;
  wire                when_MemoryEngine_l246_98;
  wire                when_MemoryEngine_l246_99;
  wire                when_MemoryEngine_l246_100;
  wire                when_MemoryEngine_l246_101;
  wire                when_MemoryEngine_l246_102;
  wire                when_MemoryEngine_l246_103;
  wire                when_MemoryEngine_l246_104;
  wire                when_MemoryEngine_l246_105;
  wire                when_MemoryEngine_l246_106;
  wire                when_MemoryEngine_l246_107;
  wire                when_MemoryEngine_l246_108;
  wire                when_MemoryEngine_l246_109;
  wire                when_MemoryEngine_l246_110;
  wire                when_MemoryEngine_l246_111;
  wire       [3:0]    _zz_when_MemoryEngine_l246_7;
  wire                when_MemoryEngine_l246_112;
  wire                when_MemoryEngine_l246_113;
  wire                when_MemoryEngine_l246_114;
  wire                when_MemoryEngine_l246_115;
  wire                when_MemoryEngine_l246_116;
  wire                when_MemoryEngine_l246_117;
  wire                when_MemoryEngine_l246_118;
  wire                when_MemoryEngine_l246_119;
  wire                when_MemoryEngine_l246_120;
  wire                when_MemoryEngine_l246_121;
  wire                when_MemoryEngine_l246_122;
  wire                when_MemoryEngine_l246_123;
  wire                when_MemoryEngine_l246_124;
  wire                when_MemoryEngine_l246_125;
  wire                when_MemoryEngine_l246_126;
  wire                when_MemoryEngine_l246_127;
  reg        [1:0]    state;
  reg        [31:0]   capStoreReq_axiAddr;
  reg        [511:0]  capStoreReq_wdata;
  reg        [63:0]   capStoreReq_wstrb;
  reg                 awAccepted;
  reg                 wAccepted;
  wire                when_MemoryEngine_l285;
  wire                when_MemoryEngine_l291;
  wire                when_MemoryEngine_l292;
  reg        [31:0]   _zz_io_loadWriteReqs_0_payload_data;
  wire                when_MemoryEngine_l297;
  wire                when_MemoryEngine_l297_1;
  wire                when_MemoryEngine_l297_2;
  wire                when_MemoryEngine_l297_3;
  wire                when_MemoryEngine_l297_4;
  wire                when_MemoryEngine_l297_5;
  wire                when_MemoryEngine_l297_6;
  wire                when_MemoryEngine_l297_7;
  wire                when_MemoryEngine_l297_8;
  wire                when_MemoryEngine_l297_9;
  wire                when_MemoryEngine_l297_10;
  wire                when_MemoryEngine_l297_11;
  wire                when_MemoryEngine_l297_12;
  wire                when_MemoryEngine_l297_13;
  wire                when_MemoryEngine_l297_14;
  wire                when_MemoryEngine_l297_15;
  reg        [31:0]   _zz_io_vloadWriteReqs_0_0_payload_data;
  wire       [3:0]    _zz_when_MemoryEngine_l311;
  wire                when_MemoryEngine_l311;
  wire                when_MemoryEngine_l311_1;
  wire                when_MemoryEngine_l311_2;
  wire                when_MemoryEngine_l311_3;
  wire                when_MemoryEngine_l311_4;
  wire                when_MemoryEngine_l311_5;
  wire                when_MemoryEngine_l311_6;
  wire                when_MemoryEngine_l311_7;
  wire                when_MemoryEngine_l311_8;
  wire                when_MemoryEngine_l311_9;
  wire                when_MemoryEngine_l311_10;
  wire                when_MemoryEngine_l311_11;
  wire                when_MemoryEngine_l311_12;
  wire                when_MemoryEngine_l311_13;
  wire                when_MemoryEngine_l311_14;
  wire                when_MemoryEngine_l311_15;
  reg        [31:0]   _zz_io_vloadWriteReqs_0_1_payload_data;
  wire       [3:0]    _zz_when_MemoryEngine_l311_1;
  wire                when_MemoryEngine_l311_16;
  wire                when_MemoryEngine_l311_17;
  wire                when_MemoryEngine_l311_18;
  wire                when_MemoryEngine_l311_19;
  wire                when_MemoryEngine_l311_20;
  wire                when_MemoryEngine_l311_21;
  wire                when_MemoryEngine_l311_22;
  wire                when_MemoryEngine_l311_23;
  wire                when_MemoryEngine_l311_24;
  wire                when_MemoryEngine_l311_25;
  wire                when_MemoryEngine_l311_26;
  wire                when_MemoryEngine_l311_27;
  wire                when_MemoryEngine_l311_28;
  wire                when_MemoryEngine_l311_29;
  wire                when_MemoryEngine_l311_30;
  wire                when_MemoryEngine_l311_31;
  reg        [31:0]   _zz_io_vloadWriteReqs_0_2_payload_data;
  wire       [3:0]    _zz_when_MemoryEngine_l311_2;
  wire                when_MemoryEngine_l311_32;
  wire                when_MemoryEngine_l311_33;
  wire                when_MemoryEngine_l311_34;
  wire                when_MemoryEngine_l311_35;
  wire                when_MemoryEngine_l311_36;
  wire                when_MemoryEngine_l311_37;
  wire                when_MemoryEngine_l311_38;
  wire                when_MemoryEngine_l311_39;
  wire                when_MemoryEngine_l311_40;
  wire                when_MemoryEngine_l311_41;
  wire                when_MemoryEngine_l311_42;
  wire                when_MemoryEngine_l311_43;
  wire                when_MemoryEngine_l311_44;
  wire                when_MemoryEngine_l311_45;
  wire                when_MemoryEngine_l311_46;
  wire                when_MemoryEngine_l311_47;
  reg        [31:0]   _zz_io_vloadWriteReqs_0_3_payload_data;
  wire       [3:0]    _zz_when_MemoryEngine_l311_3;
  wire                when_MemoryEngine_l311_48;
  wire                when_MemoryEngine_l311_49;
  wire                when_MemoryEngine_l311_50;
  wire                when_MemoryEngine_l311_51;
  wire                when_MemoryEngine_l311_52;
  wire                when_MemoryEngine_l311_53;
  wire                when_MemoryEngine_l311_54;
  wire                when_MemoryEngine_l311_55;
  wire                when_MemoryEngine_l311_56;
  wire                when_MemoryEngine_l311_57;
  wire                when_MemoryEngine_l311_58;
  wire                when_MemoryEngine_l311_59;
  wire                when_MemoryEngine_l311_60;
  wire                when_MemoryEngine_l311_61;
  wire                when_MemoryEngine_l311_62;
  wire                when_MemoryEngine_l311_63;
  reg        [31:0]   _zz_io_vloadWriteReqs_0_4_payload_data;
  wire       [3:0]    _zz_when_MemoryEngine_l311_4;
  wire                when_MemoryEngine_l311_64;
  wire                when_MemoryEngine_l311_65;
  wire                when_MemoryEngine_l311_66;
  wire                when_MemoryEngine_l311_67;
  wire                when_MemoryEngine_l311_68;
  wire                when_MemoryEngine_l311_69;
  wire                when_MemoryEngine_l311_70;
  wire                when_MemoryEngine_l311_71;
  wire                when_MemoryEngine_l311_72;
  wire                when_MemoryEngine_l311_73;
  wire                when_MemoryEngine_l311_74;
  wire                when_MemoryEngine_l311_75;
  wire                when_MemoryEngine_l311_76;
  wire                when_MemoryEngine_l311_77;
  wire                when_MemoryEngine_l311_78;
  wire                when_MemoryEngine_l311_79;
  reg        [31:0]   _zz_io_vloadWriteReqs_0_5_payload_data;
  wire       [3:0]    _zz_when_MemoryEngine_l311_5;
  wire                when_MemoryEngine_l311_80;
  wire                when_MemoryEngine_l311_81;
  wire                when_MemoryEngine_l311_82;
  wire                when_MemoryEngine_l311_83;
  wire                when_MemoryEngine_l311_84;
  wire                when_MemoryEngine_l311_85;
  wire                when_MemoryEngine_l311_86;
  wire                when_MemoryEngine_l311_87;
  wire                when_MemoryEngine_l311_88;
  wire                when_MemoryEngine_l311_89;
  wire                when_MemoryEngine_l311_90;
  wire                when_MemoryEngine_l311_91;
  wire                when_MemoryEngine_l311_92;
  wire                when_MemoryEngine_l311_93;
  wire                when_MemoryEngine_l311_94;
  wire                when_MemoryEngine_l311_95;
  reg        [31:0]   _zz_io_vloadWriteReqs_0_6_payload_data;
  wire       [3:0]    _zz_when_MemoryEngine_l311_6;
  wire                when_MemoryEngine_l311_96;
  wire                when_MemoryEngine_l311_97;
  wire                when_MemoryEngine_l311_98;
  wire                when_MemoryEngine_l311_99;
  wire                when_MemoryEngine_l311_100;
  wire                when_MemoryEngine_l311_101;
  wire                when_MemoryEngine_l311_102;
  wire                when_MemoryEngine_l311_103;
  wire                when_MemoryEngine_l311_104;
  wire                when_MemoryEngine_l311_105;
  wire                when_MemoryEngine_l311_106;
  wire                when_MemoryEngine_l311_107;
  wire                when_MemoryEngine_l311_108;
  wire                when_MemoryEngine_l311_109;
  wire                when_MemoryEngine_l311_110;
  wire                when_MemoryEngine_l311_111;
  reg        [31:0]   _zz_io_vloadWriteReqs_0_7_payload_data;
  wire       [3:0]    _zz_when_MemoryEngine_l311_7;
  wire                when_MemoryEngine_l311_112;
  wire                when_MemoryEngine_l311_113;
  wire                when_MemoryEngine_l311_114;
  wire                when_MemoryEngine_l311_115;
  wire                when_MemoryEngine_l311_116;
  wire                when_MemoryEngine_l311_117;
  wire                when_MemoryEngine_l311_118;
  wire                when_MemoryEngine_l311_119;
  wire                when_MemoryEngine_l311_120;
  wire                when_MemoryEngine_l311_121;
  wire                when_MemoryEngine_l311_122;
  wire                when_MemoryEngine_l311_123;
  wire                when_MemoryEngine_l311_124;
  wire                when_MemoryEngine_l311_125;
  wire                when_MemoryEngine_l311_126;
  wire                when_MemoryEngine_l311_127;
  wire                when_MemoryEngine_l340;
  wire                when_MemoryEngine_l341;
  wire                io_axiMaster_aw_fire;
  wire                io_axiMaster_w_fire;
  wire                when_MemoryEngine_l353;
  `ifndef SYNTHESIS
  reg [79:0] state_string;
  `endif


  assign _zz__zz_loadReqEntry_wordOff = ({2'd0,io_loadAddrData_0} <<< 2'd2);
  assign _zz_loadReqEntry_wordOff_1 = (_zz_loadReqEntry_wordOff >>> 2'd2);
  assign _zz__zz_loadReqEntry_axiAddr_2 = ({2'd0,_zz__zz_loadReqEntry_axiAddr_2_1} <<< 2'd2);
  assign _zz__zz_loadReqEntry_axiAddr_2_1 = (io_loadAddrData_0 + _zz__zz_loadReqEntry_axiAddr_2_2);
  assign _zz__zz_loadReqEntry_axiAddr_2_2 = {29'd0, io_loadSlots_0_offset};
  assign _zz_loadReqEntry_destAddr = {8'd0, io_loadSlots_0_offset};
  assign _zz_loadReqEntry_wordOff_2 = (_zz_loadReqEntry_axiAddr_2 >>> 2'd2);
  assign _zz__zz_io_push_payload_axiAddr_1 = ({2'd0,io_storeAddrData_0} <<< 2'd2);
  assign _zz__zz_when_MemoryEngine_l235 = (_zz_io_push_payload_axiAddr_1 >>> 2'd2);
  StreamFifo storeReqFifo (
    .io_push_valid           (storeReqFifo_io_push_valid                ), //i
    .io_push_ready           (storeReqFifo_io_push_ready                ), //o
    .io_push_payload_axiAddr (storeReqFifo_io_push_payload_axiAddr[31:0]), //i
    .io_push_payload_wdata   (storeReqFifo_io_push_payload_wdata[511:0] ), //i
    .io_push_payload_wstrb   (storeReqFifo_io_push_payload_wstrb[63:0]  ), //i
    .io_pop_valid            (storeReqFifo_io_pop_valid                 ), //o
    .io_pop_ready            (storeReqFifo_io_pop_ready                 ), //i
    .io_pop_payload_axiAddr  (storeReqFifo_io_pop_payload_axiAddr[31:0] ), //o
    .io_pop_payload_wdata    (storeReqFifo_io_pop_payload_wdata[511:0]  ), //o
    .io_pop_payload_wstrb    (storeReqFifo_io_pop_payload_wstrb[63:0]   ), //o
    .io_flush                (1'b0                                      ), //i
    .io_occupancy            (storeReqFifo_io_occupancy[3:0]            ), //o
    .io_availability         (storeReqFifo_io_availability[3:0]         ), //o
    .clk                     (clk                                       ), //i
    .reset                   (reset                                     )  //i
  );
  `ifndef SYNTHESIS
  always @(*) begin
    case(state)
      MemState_IDLE : state_string = "IDLE      ";
      MemState_STORE_AW_W : state_string = "STORE_AW_W";
      MemState_STORE_B : state_string = "STORE_B   ";
      default : state_string = "??????????";
    endcase
  end
  `endif

  assign axiSizeVal = 3'b110;
  always @(*) begin
    io_stall = 1'b0;
    if(when_MemoryEngine_l167) begin
      io_stall = 1'b1;
    end
    if(when_MemoryEngine_l172) begin
      io_stall = 1'b1;
    end
  end

  always @(*) begin
    io_loadWriteReqs_0_valid = 1'b0;
    if(when_MemoryEngine_l285) begin
      if(when_MemoryEngine_l291) begin
        if(when_MemoryEngine_l292) begin
          io_loadWriteReqs_0_valid = 1'b1;
        end
      end
    end
  end

  always @(*) begin
    io_loadWriteReqs_0_payload_addr = 11'h0;
    if(when_MemoryEngine_l285) begin
      if(when_MemoryEngine_l291) begin
        if(when_MemoryEngine_l292) begin
          io_loadWriteReqs_0_payload_addr = loadReqEntry_destAddr;
        end
      end
    end
  end

  always @(*) begin
    io_loadWriteReqs_0_payload_data = 32'h0;
    if(when_MemoryEngine_l285) begin
      if(when_MemoryEngine_l291) begin
        if(when_MemoryEngine_l292) begin
          io_loadWriteReqs_0_payload_data = _zz_io_loadWriteReqs_0_payload_data;
        end
      end
    end
  end

  always @(*) begin
    io_constWriteReqs_0_valid = 1'b0;
    if(when_MemoryEngine_l103) begin
      io_constWriteReqs_0_valid = 1'b1;
    end
  end

  always @(*) begin
    io_constWriteReqs_0_payload_addr = 11'h0;
    if(when_MemoryEngine_l103) begin
      io_constWriteReqs_0_payload_addr = io_loadSlots_0_dest;
    end
  end

  always @(*) begin
    io_constWriteReqs_0_payload_data = 32'h0;
    if(when_MemoryEngine_l103) begin
      io_constWriteReqs_0_payload_data = io_loadSlots_0_immediate;
    end
  end

  always @(*) begin
    io_vloadWriteReqs_0_0_valid = 1'b0;
    if(when_MemoryEngine_l285) begin
      if(when_MemoryEngine_l291) begin
        if(!when_MemoryEngine_l292) begin
          io_vloadWriteReqs_0_0_valid = 1'b1;
        end
      end
    end
  end

  always @(*) begin
    io_vloadWriteReqs_0_0_payload_addr = 11'h0;
    if(when_MemoryEngine_l285) begin
      if(when_MemoryEngine_l291) begin
        if(!when_MemoryEngine_l292) begin
          io_vloadWriteReqs_0_0_payload_addr = (loadReqEntry_destAddr + 11'h0);
        end
      end
    end
  end

  always @(*) begin
    io_vloadWriteReqs_0_0_payload_data = 32'h0;
    if(when_MemoryEngine_l285) begin
      if(when_MemoryEngine_l291) begin
        if(!when_MemoryEngine_l292) begin
          io_vloadWriteReqs_0_0_payload_data = _zz_io_vloadWriteReqs_0_0_payload_data;
        end
      end
    end
  end

  always @(*) begin
    io_vloadWriteReqs_0_1_valid = 1'b0;
    if(when_MemoryEngine_l285) begin
      if(when_MemoryEngine_l291) begin
        if(!when_MemoryEngine_l292) begin
          io_vloadWriteReqs_0_1_valid = 1'b1;
        end
      end
    end
  end

  always @(*) begin
    io_vloadWriteReqs_0_1_payload_addr = 11'h0;
    if(when_MemoryEngine_l285) begin
      if(when_MemoryEngine_l291) begin
        if(!when_MemoryEngine_l292) begin
          io_vloadWriteReqs_0_1_payload_addr = (loadReqEntry_destAddr + 11'h001);
        end
      end
    end
  end

  always @(*) begin
    io_vloadWriteReqs_0_1_payload_data = 32'h0;
    if(when_MemoryEngine_l285) begin
      if(when_MemoryEngine_l291) begin
        if(!when_MemoryEngine_l292) begin
          io_vloadWriteReqs_0_1_payload_data = _zz_io_vloadWriteReqs_0_1_payload_data;
        end
      end
    end
  end

  always @(*) begin
    io_vloadWriteReqs_0_2_valid = 1'b0;
    if(when_MemoryEngine_l285) begin
      if(when_MemoryEngine_l291) begin
        if(!when_MemoryEngine_l292) begin
          io_vloadWriteReqs_0_2_valid = 1'b1;
        end
      end
    end
  end

  always @(*) begin
    io_vloadWriteReqs_0_2_payload_addr = 11'h0;
    if(when_MemoryEngine_l285) begin
      if(when_MemoryEngine_l291) begin
        if(!when_MemoryEngine_l292) begin
          io_vloadWriteReqs_0_2_payload_addr = (loadReqEntry_destAddr + 11'h002);
        end
      end
    end
  end

  always @(*) begin
    io_vloadWriteReqs_0_2_payload_data = 32'h0;
    if(when_MemoryEngine_l285) begin
      if(when_MemoryEngine_l291) begin
        if(!when_MemoryEngine_l292) begin
          io_vloadWriteReqs_0_2_payload_data = _zz_io_vloadWriteReqs_0_2_payload_data;
        end
      end
    end
  end

  always @(*) begin
    io_vloadWriteReqs_0_3_valid = 1'b0;
    if(when_MemoryEngine_l285) begin
      if(when_MemoryEngine_l291) begin
        if(!when_MemoryEngine_l292) begin
          io_vloadWriteReqs_0_3_valid = 1'b1;
        end
      end
    end
  end

  always @(*) begin
    io_vloadWriteReqs_0_3_payload_addr = 11'h0;
    if(when_MemoryEngine_l285) begin
      if(when_MemoryEngine_l291) begin
        if(!when_MemoryEngine_l292) begin
          io_vloadWriteReqs_0_3_payload_addr = (loadReqEntry_destAddr + 11'h003);
        end
      end
    end
  end

  always @(*) begin
    io_vloadWriteReqs_0_3_payload_data = 32'h0;
    if(when_MemoryEngine_l285) begin
      if(when_MemoryEngine_l291) begin
        if(!when_MemoryEngine_l292) begin
          io_vloadWriteReqs_0_3_payload_data = _zz_io_vloadWriteReqs_0_3_payload_data;
        end
      end
    end
  end

  always @(*) begin
    io_vloadWriteReqs_0_4_valid = 1'b0;
    if(when_MemoryEngine_l285) begin
      if(when_MemoryEngine_l291) begin
        if(!when_MemoryEngine_l292) begin
          io_vloadWriteReqs_0_4_valid = 1'b1;
        end
      end
    end
  end

  always @(*) begin
    io_vloadWriteReqs_0_4_payload_addr = 11'h0;
    if(when_MemoryEngine_l285) begin
      if(when_MemoryEngine_l291) begin
        if(!when_MemoryEngine_l292) begin
          io_vloadWriteReqs_0_4_payload_addr = (loadReqEntry_destAddr + 11'h004);
        end
      end
    end
  end

  always @(*) begin
    io_vloadWriteReqs_0_4_payload_data = 32'h0;
    if(when_MemoryEngine_l285) begin
      if(when_MemoryEngine_l291) begin
        if(!when_MemoryEngine_l292) begin
          io_vloadWriteReqs_0_4_payload_data = _zz_io_vloadWriteReqs_0_4_payload_data;
        end
      end
    end
  end

  always @(*) begin
    io_vloadWriteReqs_0_5_valid = 1'b0;
    if(when_MemoryEngine_l285) begin
      if(when_MemoryEngine_l291) begin
        if(!when_MemoryEngine_l292) begin
          io_vloadWriteReqs_0_5_valid = 1'b1;
        end
      end
    end
  end

  always @(*) begin
    io_vloadWriteReqs_0_5_payload_addr = 11'h0;
    if(when_MemoryEngine_l285) begin
      if(when_MemoryEngine_l291) begin
        if(!when_MemoryEngine_l292) begin
          io_vloadWriteReqs_0_5_payload_addr = (loadReqEntry_destAddr + 11'h005);
        end
      end
    end
  end

  always @(*) begin
    io_vloadWriteReqs_0_5_payload_data = 32'h0;
    if(when_MemoryEngine_l285) begin
      if(when_MemoryEngine_l291) begin
        if(!when_MemoryEngine_l292) begin
          io_vloadWriteReqs_0_5_payload_data = _zz_io_vloadWriteReqs_0_5_payload_data;
        end
      end
    end
  end

  always @(*) begin
    io_vloadWriteReqs_0_6_valid = 1'b0;
    if(when_MemoryEngine_l285) begin
      if(when_MemoryEngine_l291) begin
        if(!when_MemoryEngine_l292) begin
          io_vloadWriteReqs_0_6_valid = 1'b1;
        end
      end
    end
  end

  always @(*) begin
    io_vloadWriteReqs_0_6_payload_addr = 11'h0;
    if(when_MemoryEngine_l285) begin
      if(when_MemoryEngine_l291) begin
        if(!when_MemoryEngine_l292) begin
          io_vloadWriteReqs_0_6_payload_addr = (loadReqEntry_destAddr + 11'h006);
        end
      end
    end
  end

  always @(*) begin
    io_vloadWriteReqs_0_6_payload_data = 32'h0;
    if(when_MemoryEngine_l285) begin
      if(when_MemoryEngine_l291) begin
        if(!when_MemoryEngine_l292) begin
          io_vloadWriteReqs_0_6_payload_data = _zz_io_vloadWriteReqs_0_6_payload_data;
        end
      end
    end
  end

  always @(*) begin
    io_vloadWriteReqs_0_7_valid = 1'b0;
    if(when_MemoryEngine_l285) begin
      if(when_MemoryEngine_l291) begin
        if(!when_MemoryEngine_l292) begin
          io_vloadWriteReqs_0_7_valid = 1'b1;
        end
      end
    end
  end

  always @(*) begin
    io_vloadWriteReqs_0_7_payload_addr = 11'h0;
    if(when_MemoryEngine_l285) begin
      if(when_MemoryEngine_l291) begin
        if(!when_MemoryEngine_l292) begin
          io_vloadWriteReqs_0_7_payload_addr = (loadReqEntry_destAddr + 11'h007);
        end
      end
    end
  end

  always @(*) begin
    io_vloadWriteReqs_0_7_payload_data = 32'h0;
    if(when_MemoryEngine_l285) begin
      if(when_MemoryEngine_l291) begin
        if(!when_MemoryEngine_l292) begin
          io_vloadWriteReqs_0_7_payload_data = _zz_io_vloadWriteReqs_0_7_payload_data;
        end
      end
    end
  end

  always @(*) begin
    io_axiMaster_aw_valid = 1'b0;
    case(state)
      MemState_IDLE : begin
      end
      MemState_STORE_AW_W : begin
        if(when_MemoryEngine_l340) begin
          io_axiMaster_aw_valid = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_axiMaster_aw_payload_addr = 32'h0;
    case(state)
      MemState_IDLE : begin
      end
      MemState_STORE_AW_W : begin
        io_axiMaster_aw_payload_addr = capStoreReq_axiAddr;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_axiMaster_aw_payload_len = 8'h0;
    case(state)
      MemState_IDLE : begin
      end
      MemState_STORE_AW_W : begin
        io_axiMaster_aw_payload_len = 8'h0;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_axiMaster_aw_payload_size = axiSizeVal;
    case(state)
      MemState_IDLE : begin
      end
      MemState_STORE_AW_W : begin
        io_axiMaster_aw_payload_size = axiSizeVal;
      end
      default : begin
      end
    endcase
  end

  assign io_axiMaster_aw_payload_burst = 2'b01;
  assign io_axiMaster_aw_payload_id = 4'b0000;
  always @(*) begin
    io_axiMaster_w_valid = 1'b0;
    case(state)
      MemState_IDLE : begin
      end
      MemState_STORE_AW_W : begin
        if(when_MemoryEngine_l341) begin
          io_axiMaster_w_valid = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_axiMaster_w_payload_data = 512'h0;
    case(state)
      MemState_IDLE : begin
      end
      MemState_STORE_AW_W : begin
        io_axiMaster_w_payload_data = capStoreReq_wdata;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_axiMaster_w_payload_strb = 64'h0;
    case(state)
      MemState_IDLE : begin
      end
      MemState_STORE_AW_W : begin
        io_axiMaster_w_payload_strb = capStoreReq_wstrb;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_axiMaster_w_payload_last = 1'b1;
    case(state)
      MemState_IDLE : begin
      end
      MemState_STORE_AW_W : begin
        io_axiMaster_w_payload_last = 1'b1;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_axiMaster_b_ready = 1'b0;
    case(state)
      MemState_IDLE : begin
      end
      MemState_STORE_AW_W : begin
      end
      default : begin
        io_axiMaster_b_ready = 1'b1;
      end
    endcase
  end

  assign when_MemoryEngine_l103 = ((io_loadSlots_0_valid && io_valid) && (io_loadSlots_0_opcode == 3'b100));
  always @(*) begin
    storeReqFifo_io_push_valid = 1'b0;
    if(when_MemoryEngine_l215) begin
      storeReqFifo_io_push_valid = 1'b1;
    end
  end

  assign _zz_io_push_payload_axiAddr = 608'h0;
  always @(*) begin
    storeReqFifo_io_push_payload_axiAddr = _zz_io_push_payload_axiAddr[31 : 0];
    if(when_MemoryEngine_l215) begin
      storeReqFifo_io_push_payload_axiAddr = (_zz_io_push_payload_axiAddr_1 & (~ 32'h0000003f));
    end
  end

  always @(*) begin
    storeReqFifo_io_push_payload_wdata = _zz_io_push_payload_axiAddr[543 : 32];
    if(when_MemoryEngine_l215) begin
      storeReqFifo_io_push_payload_wdata = _zz_io_push_payload_wdata;
    end
  end

  always @(*) begin
    storeReqFifo_io_push_payload_wstrb = _zz_io_push_payload_axiAddr[607 : 544];
    if(when_MemoryEngine_l215) begin
      storeReqFifo_io_push_payload_wstrb = _zz_io_push_payload_wstrb;
    end
  end

  always @(*) begin
    anyLoadOp = 1'b0;
    if(isLoadOp_0) begin
      anyLoadOp = 1'b1;
    end
  end

  assign isLoadOp_0 = ((io_loadSlots_0_valid && io_valid) && (((io_loadSlots_0_opcode == 3'b001) || (io_loadSlots_0_opcode == 3'b010)) || (io_loadSlots_0_opcode == 3'b011)));
  always @(*) begin
    anyStoreOp = 1'b0;
    if(isStoreOp_0) begin
      anyStoreOp = 1'b1;
    end
  end

  assign isStoreOp_0 = ((io_storeSlots_0_valid && io_valid) && ((io_storeSlots_0_opcode == 2'b01) || (io_storeSlots_0_opcode == 2'b10)));
  assign when_MemoryEngine_l167 = (anyLoadOp && loadReqValid);
  assign when_MemoryEngine_l172 = (anyStoreOp && (! storeReqFifo_io_push_ready));
  assign when_MemoryEngine_l180 = (isLoadOp_0 && (! io_stall));
  assign _zz_loadReqEntry_wordOff = _zz__zz_loadReqEntry_wordOff[31:0];
  assign _zz_loadReqEntry_axiAddr = 32'h0000003f;
  assign _zz_loadReqEntry_axiAddr_1 = (_zz_loadReqEntry_wordOff & (~ _zz_loadReqEntry_axiAddr));
  assign _zz_loadReqEntry_axiAddr_2 = _zz__zz_loadReqEntry_axiAddr_2[31:0];
  assign when_MemoryEngine_l215 = (isStoreOp_0 && (! io_stall));
  assign _zz_io_push_payload_axiAddr_1 = _zz__zz_io_push_payload_axiAddr_1[31:0];
  assign _zz_when_MemoryEngine_l235 = _zz__zz_when_MemoryEngine_l235[3:0];
  always @(*) begin
    _zz_io_push_payload_wdata = 512'h0;
    case(io_storeSlots_0_opcode)
      2'b01 : begin
        if(when_MemoryEngine_l235) begin
          _zz_io_push_payload_wdata[31 : 0] = io_storeSrcData_0;
        end
        if(when_MemoryEngine_l235_1) begin
          _zz_io_push_payload_wdata[63 : 32] = io_storeSrcData_0;
        end
        if(when_MemoryEngine_l235_2) begin
          _zz_io_push_payload_wdata[95 : 64] = io_storeSrcData_0;
        end
        if(when_MemoryEngine_l235_3) begin
          _zz_io_push_payload_wdata[127 : 96] = io_storeSrcData_0;
        end
        if(when_MemoryEngine_l235_4) begin
          _zz_io_push_payload_wdata[159 : 128] = io_storeSrcData_0;
        end
        if(when_MemoryEngine_l235_5) begin
          _zz_io_push_payload_wdata[191 : 160] = io_storeSrcData_0;
        end
        if(when_MemoryEngine_l235_6) begin
          _zz_io_push_payload_wdata[223 : 192] = io_storeSrcData_0;
        end
        if(when_MemoryEngine_l235_7) begin
          _zz_io_push_payload_wdata[255 : 224] = io_storeSrcData_0;
        end
        if(when_MemoryEngine_l235_8) begin
          _zz_io_push_payload_wdata[287 : 256] = io_storeSrcData_0;
        end
        if(when_MemoryEngine_l235_9) begin
          _zz_io_push_payload_wdata[319 : 288] = io_storeSrcData_0;
        end
        if(when_MemoryEngine_l235_10) begin
          _zz_io_push_payload_wdata[351 : 320] = io_storeSrcData_0;
        end
        if(when_MemoryEngine_l235_11) begin
          _zz_io_push_payload_wdata[383 : 352] = io_storeSrcData_0;
        end
        if(when_MemoryEngine_l235_12) begin
          _zz_io_push_payload_wdata[415 : 384] = io_storeSrcData_0;
        end
        if(when_MemoryEngine_l235_13) begin
          _zz_io_push_payload_wdata[447 : 416] = io_storeSrcData_0;
        end
        if(when_MemoryEngine_l235_14) begin
          _zz_io_push_payload_wdata[479 : 448] = io_storeSrcData_0;
        end
        if(when_MemoryEngine_l235_15) begin
          _zz_io_push_payload_wdata[511 : 480] = io_storeSrcData_0;
        end
      end
      2'b10 : begin
        if(when_MemoryEngine_l246) begin
          _zz_io_push_payload_wdata[31 : 0] = io_vstoreSrcData_0_0;
        end
        if(when_MemoryEngine_l246_1) begin
          _zz_io_push_payload_wdata[63 : 32] = io_vstoreSrcData_0_0;
        end
        if(when_MemoryEngine_l246_2) begin
          _zz_io_push_payload_wdata[95 : 64] = io_vstoreSrcData_0_0;
        end
        if(when_MemoryEngine_l246_3) begin
          _zz_io_push_payload_wdata[127 : 96] = io_vstoreSrcData_0_0;
        end
        if(when_MemoryEngine_l246_4) begin
          _zz_io_push_payload_wdata[159 : 128] = io_vstoreSrcData_0_0;
        end
        if(when_MemoryEngine_l246_5) begin
          _zz_io_push_payload_wdata[191 : 160] = io_vstoreSrcData_0_0;
        end
        if(when_MemoryEngine_l246_6) begin
          _zz_io_push_payload_wdata[223 : 192] = io_vstoreSrcData_0_0;
        end
        if(when_MemoryEngine_l246_7) begin
          _zz_io_push_payload_wdata[255 : 224] = io_vstoreSrcData_0_0;
        end
        if(when_MemoryEngine_l246_8) begin
          _zz_io_push_payload_wdata[287 : 256] = io_vstoreSrcData_0_0;
        end
        if(when_MemoryEngine_l246_9) begin
          _zz_io_push_payload_wdata[319 : 288] = io_vstoreSrcData_0_0;
        end
        if(when_MemoryEngine_l246_10) begin
          _zz_io_push_payload_wdata[351 : 320] = io_vstoreSrcData_0_0;
        end
        if(when_MemoryEngine_l246_11) begin
          _zz_io_push_payload_wdata[383 : 352] = io_vstoreSrcData_0_0;
        end
        if(when_MemoryEngine_l246_12) begin
          _zz_io_push_payload_wdata[415 : 384] = io_vstoreSrcData_0_0;
        end
        if(when_MemoryEngine_l246_13) begin
          _zz_io_push_payload_wdata[447 : 416] = io_vstoreSrcData_0_0;
        end
        if(when_MemoryEngine_l246_14) begin
          _zz_io_push_payload_wdata[479 : 448] = io_vstoreSrcData_0_0;
        end
        if(when_MemoryEngine_l246_15) begin
          _zz_io_push_payload_wdata[511 : 480] = io_vstoreSrcData_0_0;
        end
        if(when_MemoryEngine_l246_16) begin
          _zz_io_push_payload_wdata[31 : 0] = io_vstoreSrcData_0_1;
        end
        if(when_MemoryEngine_l246_17) begin
          _zz_io_push_payload_wdata[63 : 32] = io_vstoreSrcData_0_1;
        end
        if(when_MemoryEngine_l246_18) begin
          _zz_io_push_payload_wdata[95 : 64] = io_vstoreSrcData_0_1;
        end
        if(when_MemoryEngine_l246_19) begin
          _zz_io_push_payload_wdata[127 : 96] = io_vstoreSrcData_0_1;
        end
        if(when_MemoryEngine_l246_20) begin
          _zz_io_push_payload_wdata[159 : 128] = io_vstoreSrcData_0_1;
        end
        if(when_MemoryEngine_l246_21) begin
          _zz_io_push_payload_wdata[191 : 160] = io_vstoreSrcData_0_1;
        end
        if(when_MemoryEngine_l246_22) begin
          _zz_io_push_payload_wdata[223 : 192] = io_vstoreSrcData_0_1;
        end
        if(when_MemoryEngine_l246_23) begin
          _zz_io_push_payload_wdata[255 : 224] = io_vstoreSrcData_0_1;
        end
        if(when_MemoryEngine_l246_24) begin
          _zz_io_push_payload_wdata[287 : 256] = io_vstoreSrcData_0_1;
        end
        if(when_MemoryEngine_l246_25) begin
          _zz_io_push_payload_wdata[319 : 288] = io_vstoreSrcData_0_1;
        end
        if(when_MemoryEngine_l246_26) begin
          _zz_io_push_payload_wdata[351 : 320] = io_vstoreSrcData_0_1;
        end
        if(when_MemoryEngine_l246_27) begin
          _zz_io_push_payload_wdata[383 : 352] = io_vstoreSrcData_0_1;
        end
        if(when_MemoryEngine_l246_28) begin
          _zz_io_push_payload_wdata[415 : 384] = io_vstoreSrcData_0_1;
        end
        if(when_MemoryEngine_l246_29) begin
          _zz_io_push_payload_wdata[447 : 416] = io_vstoreSrcData_0_1;
        end
        if(when_MemoryEngine_l246_30) begin
          _zz_io_push_payload_wdata[479 : 448] = io_vstoreSrcData_0_1;
        end
        if(when_MemoryEngine_l246_31) begin
          _zz_io_push_payload_wdata[511 : 480] = io_vstoreSrcData_0_1;
        end
        if(when_MemoryEngine_l246_32) begin
          _zz_io_push_payload_wdata[31 : 0] = io_vstoreSrcData_0_2;
        end
        if(when_MemoryEngine_l246_33) begin
          _zz_io_push_payload_wdata[63 : 32] = io_vstoreSrcData_0_2;
        end
        if(when_MemoryEngine_l246_34) begin
          _zz_io_push_payload_wdata[95 : 64] = io_vstoreSrcData_0_2;
        end
        if(when_MemoryEngine_l246_35) begin
          _zz_io_push_payload_wdata[127 : 96] = io_vstoreSrcData_0_2;
        end
        if(when_MemoryEngine_l246_36) begin
          _zz_io_push_payload_wdata[159 : 128] = io_vstoreSrcData_0_2;
        end
        if(when_MemoryEngine_l246_37) begin
          _zz_io_push_payload_wdata[191 : 160] = io_vstoreSrcData_0_2;
        end
        if(when_MemoryEngine_l246_38) begin
          _zz_io_push_payload_wdata[223 : 192] = io_vstoreSrcData_0_2;
        end
        if(when_MemoryEngine_l246_39) begin
          _zz_io_push_payload_wdata[255 : 224] = io_vstoreSrcData_0_2;
        end
        if(when_MemoryEngine_l246_40) begin
          _zz_io_push_payload_wdata[287 : 256] = io_vstoreSrcData_0_2;
        end
        if(when_MemoryEngine_l246_41) begin
          _zz_io_push_payload_wdata[319 : 288] = io_vstoreSrcData_0_2;
        end
        if(when_MemoryEngine_l246_42) begin
          _zz_io_push_payload_wdata[351 : 320] = io_vstoreSrcData_0_2;
        end
        if(when_MemoryEngine_l246_43) begin
          _zz_io_push_payload_wdata[383 : 352] = io_vstoreSrcData_0_2;
        end
        if(when_MemoryEngine_l246_44) begin
          _zz_io_push_payload_wdata[415 : 384] = io_vstoreSrcData_0_2;
        end
        if(when_MemoryEngine_l246_45) begin
          _zz_io_push_payload_wdata[447 : 416] = io_vstoreSrcData_0_2;
        end
        if(when_MemoryEngine_l246_46) begin
          _zz_io_push_payload_wdata[479 : 448] = io_vstoreSrcData_0_2;
        end
        if(when_MemoryEngine_l246_47) begin
          _zz_io_push_payload_wdata[511 : 480] = io_vstoreSrcData_0_2;
        end
        if(when_MemoryEngine_l246_48) begin
          _zz_io_push_payload_wdata[31 : 0] = io_vstoreSrcData_0_3;
        end
        if(when_MemoryEngine_l246_49) begin
          _zz_io_push_payload_wdata[63 : 32] = io_vstoreSrcData_0_3;
        end
        if(when_MemoryEngine_l246_50) begin
          _zz_io_push_payload_wdata[95 : 64] = io_vstoreSrcData_0_3;
        end
        if(when_MemoryEngine_l246_51) begin
          _zz_io_push_payload_wdata[127 : 96] = io_vstoreSrcData_0_3;
        end
        if(when_MemoryEngine_l246_52) begin
          _zz_io_push_payload_wdata[159 : 128] = io_vstoreSrcData_0_3;
        end
        if(when_MemoryEngine_l246_53) begin
          _zz_io_push_payload_wdata[191 : 160] = io_vstoreSrcData_0_3;
        end
        if(when_MemoryEngine_l246_54) begin
          _zz_io_push_payload_wdata[223 : 192] = io_vstoreSrcData_0_3;
        end
        if(when_MemoryEngine_l246_55) begin
          _zz_io_push_payload_wdata[255 : 224] = io_vstoreSrcData_0_3;
        end
        if(when_MemoryEngine_l246_56) begin
          _zz_io_push_payload_wdata[287 : 256] = io_vstoreSrcData_0_3;
        end
        if(when_MemoryEngine_l246_57) begin
          _zz_io_push_payload_wdata[319 : 288] = io_vstoreSrcData_0_3;
        end
        if(when_MemoryEngine_l246_58) begin
          _zz_io_push_payload_wdata[351 : 320] = io_vstoreSrcData_0_3;
        end
        if(when_MemoryEngine_l246_59) begin
          _zz_io_push_payload_wdata[383 : 352] = io_vstoreSrcData_0_3;
        end
        if(when_MemoryEngine_l246_60) begin
          _zz_io_push_payload_wdata[415 : 384] = io_vstoreSrcData_0_3;
        end
        if(when_MemoryEngine_l246_61) begin
          _zz_io_push_payload_wdata[447 : 416] = io_vstoreSrcData_0_3;
        end
        if(when_MemoryEngine_l246_62) begin
          _zz_io_push_payload_wdata[479 : 448] = io_vstoreSrcData_0_3;
        end
        if(when_MemoryEngine_l246_63) begin
          _zz_io_push_payload_wdata[511 : 480] = io_vstoreSrcData_0_3;
        end
        if(when_MemoryEngine_l246_64) begin
          _zz_io_push_payload_wdata[31 : 0] = io_vstoreSrcData_0_4;
        end
        if(when_MemoryEngine_l246_65) begin
          _zz_io_push_payload_wdata[63 : 32] = io_vstoreSrcData_0_4;
        end
        if(when_MemoryEngine_l246_66) begin
          _zz_io_push_payload_wdata[95 : 64] = io_vstoreSrcData_0_4;
        end
        if(when_MemoryEngine_l246_67) begin
          _zz_io_push_payload_wdata[127 : 96] = io_vstoreSrcData_0_4;
        end
        if(when_MemoryEngine_l246_68) begin
          _zz_io_push_payload_wdata[159 : 128] = io_vstoreSrcData_0_4;
        end
        if(when_MemoryEngine_l246_69) begin
          _zz_io_push_payload_wdata[191 : 160] = io_vstoreSrcData_0_4;
        end
        if(when_MemoryEngine_l246_70) begin
          _zz_io_push_payload_wdata[223 : 192] = io_vstoreSrcData_0_4;
        end
        if(when_MemoryEngine_l246_71) begin
          _zz_io_push_payload_wdata[255 : 224] = io_vstoreSrcData_0_4;
        end
        if(when_MemoryEngine_l246_72) begin
          _zz_io_push_payload_wdata[287 : 256] = io_vstoreSrcData_0_4;
        end
        if(when_MemoryEngine_l246_73) begin
          _zz_io_push_payload_wdata[319 : 288] = io_vstoreSrcData_0_4;
        end
        if(when_MemoryEngine_l246_74) begin
          _zz_io_push_payload_wdata[351 : 320] = io_vstoreSrcData_0_4;
        end
        if(when_MemoryEngine_l246_75) begin
          _zz_io_push_payload_wdata[383 : 352] = io_vstoreSrcData_0_4;
        end
        if(when_MemoryEngine_l246_76) begin
          _zz_io_push_payload_wdata[415 : 384] = io_vstoreSrcData_0_4;
        end
        if(when_MemoryEngine_l246_77) begin
          _zz_io_push_payload_wdata[447 : 416] = io_vstoreSrcData_0_4;
        end
        if(when_MemoryEngine_l246_78) begin
          _zz_io_push_payload_wdata[479 : 448] = io_vstoreSrcData_0_4;
        end
        if(when_MemoryEngine_l246_79) begin
          _zz_io_push_payload_wdata[511 : 480] = io_vstoreSrcData_0_4;
        end
        if(when_MemoryEngine_l246_80) begin
          _zz_io_push_payload_wdata[31 : 0] = io_vstoreSrcData_0_5;
        end
        if(when_MemoryEngine_l246_81) begin
          _zz_io_push_payload_wdata[63 : 32] = io_vstoreSrcData_0_5;
        end
        if(when_MemoryEngine_l246_82) begin
          _zz_io_push_payload_wdata[95 : 64] = io_vstoreSrcData_0_5;
        end
        if(when_MemoryEngine_l246_83) begin
          _zz_io_push_payload_wdata[127 : 96] = io_vstoreSrcData_0_5;
        end
        if(when_MemoryEngine_l246_84) begin
          _zz_io_push_payload_wdata[159 : 128] = io_vstoreSrcData_0_5;
        end
        if(when_MemoryEngine_l246_85) begin
          _zz_io_push_payload_wdata[191 : 160] = io_vstoreSrcData_0_5;
        end
        if(when_MemoryEngine_l246_86) begin
          _zz_io_push_payload_wdata[223 : 192] = io_vstoreSrcData_0_5;
        end
        if(when_MemoryEngine_l246_87) begin
          _zz_io_push_payload_wdata[255 : 224] = io_vstoreSrcData_0_5;
        end
        if(when_MemoryEngine_l246_88) begin
          _zz_io_push_payload_wdata[287 : 256] = io_vstoreSrcData_0_5;
        end
        if(when_MemoryEngine_l246_89) begin
          _zz_io_push_payload_wdata[319 : 288] = io_vstoreSrcData_0_5;
        end
        if(when_MemoryEngine_l246_90) begin
          _zz_io_push_payload_wdata[351 : 320] = io_vstoreSrcData_0_5;
        end
        if(when_MemoryEngine_l246_91) begin
          _zz_io_push_payload_wdata[383 : 352] = io_vstoreSrcData_0_5;
        end
        if(when_MemoryEngine_l246_92) begin
          _zz_io_push_payload_wdata[415 : 384] = io_vstoreSrcData_0_5;
        end
        if(when_MemoryEngine_l246_93) begin
          _zz_io_push_payload_wdata[447 : 416] = io_vstoreSrcData_0_5;
        end
        if(when_MemoryEngine_l246_94) begin
          _zz_io_push_payload_wdata[479 : 448] = io_vstoreSrcData_0_5;
        end
        if(when_MemoryEngine_l246_95) begin
          _zz_io_push_payload_wdata[511 : 480] = io_vstoreSrcData_0_5;
        end
        if(when_MemoryEngine_l246_96) begin
          _zz_io_push_payload_wdata[31 : 0] = io_vstoreSrcData_0_6;
        end
        if(when_MemoryEngine_l246_97) begin
          _zz_io_push_payload_wdata[63 : 32] = io_vstoreSrcData_0_6;
        end
        if(when_MemoryEngine_l246_98) begin
          _zz_io_push_payload_wdata[95 : 64] = io_vstoreSrcData_0_6;
        end
        if(when_MemoryEngine_l246_99) begin
          _zz_io_push_payload_wdata[127 : 96] = io_vstoreSrcData_0_6;
        end
        if(when_MemoryEngine_l246_100) begin
          _zz_io_push_payload_wdata[159 : 128] = io_vstoreSrcData_0_6;
        end
        if(when_MemoryEngine_l246_101) begin
          _zz_io_push_payload_wdata[191 : 160] = io_vstoreSrcData_0_6;
        end
        if(when_MemoryEngine_l246_102) begin
          _zz_io_push_payload_wdata[223 : 192] = io_vstoreSrcData_0_6;
        end
        if(when_MemoryEngine_l246_103) begin
          _zz_io_push_payload_wdata[255 : 224] = io_vstoreSrcData_0_6;
        end
        if(when_MemoryEngine_l246_104) begin
          _zz_io_push_payload_wdata[287 : 256] = io_vstoreSrcData_0_6;
        end
        if(when_MemoryEngine_l246_105) begin
          _zz_io_push_payload_wdata[319 : 288] = io_vstoreSrcData_0_6;
        end
        if(when_MemoryEngine_l246_106) begin
          _zz_io_push_payload_wdata[351 : 320] = io_vstoreSrcData_0_6;
        end
        if(when_MemoryEngine_l246_107) begin
          _zz_io_push_payload_wdata[383 : 352] = io_vstoreSrcData_0_6;
        end
        if(when_MemoryEngine_l246_108) begin
          _zz_io_push_payload_wdata[415 : 384] = io_vstoreSrcData_0_6;
        end
        if(when_MemoryEngine_l246_109) begin
          _zz_io_push_payload_wdata[447 : 416] = io_vstoreSrcData_0_6;
        end
        if(when_MemoryEngine_l246_110) begin
          _zz_io_push_payload_wdata[479 : 448] = io_vstoreSrcData_0_6;
        end
        if(when_MemoryEngine_l246_111) begin
          _zz_io_push_payload_wdata[511 : 480] = io_vstoreSrcData_0_6;
        end
        if(when_MemoryEngine_l246_112) begin
          _zz_io_push_payload_wdata[31 : 0] = io_vstoreSrcData_0_7;
        end
        if(when_MemoryEngine_l246_113) begin
          _zz_io_push_payload_wdata[63 : 32] = io_vstoreSrcData_0_7;
        end
        if(when_MemoryEngine_l246_114) begin
          _zz_io_push_payload_wdata[95 : 64] = io_vstoreSrcData_0_7;
        end
        if(when_MemoryEngine_l246_115) begin
          _zz_io_push_payload_wdata[127 : 96] = io_vstoreSrcData_0_7;
        end
        if(when_MemoryEngine_l246_116) begin
          _zz_io_push_payload_wdata[159 : 128] = io_vstoreSrcData_0_7;
        end
        if(when_MemoryEngine_l246_117) begin
          _zz_io_push_payload_wdata[191 : 160] = io_vstoreSrcData_0_7;
        end
        if(when_MemoryEngine_l246_118) begin
          _zz_io_push_payload_wdata[223 : 192] = io_vstoreSrcData_0_7;
        end
        if(when_MemoryEngine_l246_119) begin
          _zz_io_push_payload_wdata[255 : 224] = io_vstoreSrcData_0_7;
        end
        if(when_MemoryEngine_l246_120) begin
          _zz_io_push_payload_wdata[287 : 256] = io_vstoreSrcData_0_7;
        end
        if(when_MemoryEngine_l246_121) begin
          _zz_io_push_payload_wdata[319 : 288] = io_vstoreSrcData_0_7;
        end
        if(when_MemoryEngine_l246_122) begin
          _zz_io_push_payload_wdata[351 : 320] = io_vstoreSrcData_0_7;
        end
        if(when_MemoryEngine_l246_123) begin
          _zz_io_push_payload_wdata[383 : 352] = io_vstoreSrcData_0_7;
        end
        if(when_MemoryEngine_l246_124) begin
          _zz_io_push_payload_wdata[415 : 384] = io_vstoreSrcData_0_7;
        end
        if(when_MemoryEngine_l246_125) begin
          _zz_io_push_payload_wdata[447 : 416] = io_vstoreSrcData_0_7;
        end
        if(when_MemoryEngine_l246_126) begin
          _zz_io_push_payload_wdata[479 : 448] = io_vstoreSrcData_0_7;
        end
        if(when_MemoryEngine_l246_127) begin
          _zz_io_push_payload_wdata[511 : 480] = io_vstoreSrcData_0_7;
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    _zz_io_push_payload_wstrb = 64'h0;
    case(io_storeSlots_0_opcode)
      2'b01 : begin
        if(when_MemoryEngine_l235) begin
          _zz_io_push_payload_wstrb[3 : 0] = 4'b1111;
        end
        if(when_MemoryEngine_l235_1) begin
          _zz_io_push_payload_wstrb[7 : 4] = 4'b1111;
        end
        if(when_MemoryEngine_l235_2) begin
          _zz_io_push_payload_wstrb[11 : 8] = 4'b1111;
        end
        if(when_MemoryEngine_l235_3) begin
          _zz_io_push_payload_wstrb[15 : 12] = 4'b1111;
        end
        if(when_MemoryEngine_l235_4) begin
          _zz_io_push_payload_wstrb[19 : 16] = 4'b1111;
        end
        if(when_MemoryEngine_l235_5) begin
          _zz_io_push_payload_wstrb[23 : 20] = 4'b1111;
        end
        if(when_MemoryEngine_l235_6) begin
          _zz_io_push_payload_wstrb[27 : 24] = 4'b1111;
        end
        if(when_MemoryEngine_l235_7) begin
          _zz_io_push_payload_wstrb[31 : 28] = 4'b1111;
        end
        if(when_MemoryEngine_l235_8) begin
          _zz_io_push_payload_wstrb[35 : 32] = 4'b1111;
        end
        if(when_MemoryEngine_l235_9) begin
          _zz_io_push_payload_wstrb[39 : 36] = 4'b1111;
        end
        if(when_MemoryEngine_l235_10) begin
          _zz_io_push_payload_wstrb[43 : 40] = 4'b1111;
        end
        if(when_MemoryEngine_l235_11) begin
          _zz_io_push_payload_wstrb[47 : 44] = 4'b1111;
        end
        if(when_MemoryEngine_l235_12) begin
          _zz_io_push_payload_wstrb[51 : 48] = 4'b1111;
        end
        if(when_MemoryEngine_l235_13) begin
          _zz_io_push_payload_wstrb[55 : 52] = 4'b1111;
        end
        if(when_MemoryEngine_l235_14) begin
          _zz_io_push_payload_wstrb[59 : 56] = 4'b1111;
        end
        if(when_MemoryEngine_l235_15) begin
          _zz_io_push_payload_wstrb[63 : 60] = 4'b1111;
        end
      end
      2'b10 : begin
        if(when_MemoryEngine_l246) begin
          _zz_io_push_payload_wstrb[3 : 0] = 4'b1111;
        end
        if(when_MemoryEngine_l246_1) begin
          _zz_io_push_payload_wstrb[7 : 4] = 4'b1111;
        end
        if(when_MemoryEngine_l246_2) begin
          _zz_io_push_payload_wstrb[11 : 8] = 4'b1111;
        end
        if(when_MemoryEngine_l246_3) begin
          _zz_io_push_payload_wstrb[15 : 12] = 4'b1111;
        end
        if(when_MemoryEngine_l246_4) begin
          _zz_io_push_payload_wstrb[19 : 16] = 4'b1111;
        end
        if(when_MemoryEngine_l246_5) begin
          _zz_io_push_payload_wstrb[23 : 20] = 4'b1111;
        end
        if(when_MemoryEngine_l246_6) begin
          _zz_io_push_payload_wstrb[27 : 24] = 4'b1111;
        end
        if(when_MemoryEngine_l246_7) begin
          _zz_io_push_payload_wstrb[31 : 28] = 4'b1111;
        end
        if(when_MemoryEngine_l246_8) begin
          _zz_io_push_payload_wstrb[35 : 32] = 4'b1111;
        end
        if(when_MemoryEngine_l246_9) begin
          _zz_io_push_payload_wstrb[39 : 36] = 4'b1111;
        end
        if(when_MemoryEngine_l246_10) begin
          _zz_io_push_payload_wstrb[43 : 40] = 4'b1111;
        end
        if(when_MemoryEngine_l246_11) begin
          _zz_io_push_payload_wstrb[47 : 44] = 4'b1111;
        end
        if(when_MemoryEngine_l246_12) begin
          _zz_io_push_payload_wstrb[51 : 48] = 4'b1111;
        end
        if(when_MemoryEngine_l246_13) begin
          _zz_io_push_payload_wstrb[55 : 52] = 4'b1111;
        end
        if(when_MemoryEngine_l246_14) begin
          _zz_io_push_payload_wstrb[59 : 56] = 4'b1111;
        end
        if(when_MemoryEngine_l246_15) begin
          _zz_io_push_payload_wstrb[63 : 60] = 4'b1111;
        end
        if(when_MemoryEngine_l246_16) begin
          _zz_io_push_payload_wstrb[3 : 0] = 4'b1111;
        end
        if(when_MemoryEngine_l246_17) begin
          _zz_io_push_payload_wstrb[7 : 4] = 4'b1111;
        end
        if(when_MemoryEngine_l246_18) begin
          _zz_io_push_payload_wstrb[11 : 8] = 4'b1111;
        end
        if(when_MemoryEngine_l246_19) begin
          _zz_io_push_payload_wstrb[15 : 12] = 4'b1111;
        end
        if(when_MemoryEngine_l246_20) begin
          _zz_io_push_payload_wstrb[19 : 16] = 4'b1111;
        end
        if(when_MemoryEngine_l246_21) begin
          _zz_io_push_payload_wstrb[23 : 20] = 4'b1111;
        end
        if(when_MemoryEngine_l246_22) begin
          _zz_io_push_payload_wstrb[27 : 24] = 4'b1111;
        end
        if(when_MemoryEngine_l246_23) begin
          _zz_io_push_payload_wstrb[31 : 28] = 4'b1111;
        end
        if(when_MemoryEngine_l246_24) begin
          _zz_io_push_payload_wstrb[35 : 32] = 4'b1111;
        end
        if(when_MemoryEngine_l246_25) begin
          _zz_io_push_payload_wstrb[39 : 36] = 4'b1111;
        end
        if(when_MemoryEngine_l246_26) begin
          _zz_io_push_payload_wstrb[43 : 40] = 4'b1111;
        end
        if(when_MemoryEngine_l246_27) begin
          _zz_io_push_payload_wstrb[47 : 44] = 4'b1111;
        end
        if(when_MemoryEngine_l246_28) begin
          _zz_io_push_payload_wstrb[51 : 48] = 4'b1111;
        end
        if(when_MemoryEngine_l246_29) begin
          _zz_io_push_payload_wstrb[55 : 52] = 4'b1111;
        end
        if(when_MemoryEngine_l246_30) begin
          _zz_io_push_payload_wstrb[59 : 56] = 4'b1111;
        end
        if(when_MemoryEngine_l246_31) begin
          _zz_io_push_payload_wstrb[63 : 60] = 4'b1111;
        end
        if(when_MemoryEngine_l246_32) begin
          _zz_io_push_payload_wstrb[3 : 0] = 4'b1111;
        end
        if(when_MemoryEngine_l246_33) begin
          _zz_io_push_payload_wstrb[7 : 4] = 4'b1111;
        end
        if(when_MemoryEngine_l246_34) begin
          _zz_io_push_payload_wstrb[11 : 8] = 4'b1111;
        end
        if(when_MemoryEngine_l246_35) begin
          _zz_io_push_payload_wstrb[15 : 12] = 4'b1111;
        end
        if(when_MemoryEngine_l246_36) begin
          _zz_io_push_payload_wstrb[19 : 16] = 4'b1111;
        end
        if(when_MemoryEngine_l246_37) begin
          _zz_io_push_payload_wstrb[23 : 20] = 4'b1111;
        end
        if(when_MemoryEngine_l246_38) begin
          _zz_io_push_payload_wstrb[27 : 24] = 4'b1111;
        end
        if(when_MemoryEngine_l246_39) begin
          _zz_io_push_payload_wstrb[31 : 28] = 4'b1111;
        end
        if(when_MemoryEngine_l246_40) begin
          _zz_io_push_payload_wstrb[35 : 32] = 4'b1111;
        end
        if(when_MemoryEngine_l246_41) begin
          _zz_io_push_payload_wstrb[39 : 36] = 4'b1111;
        end
        if(when_MemoryEngine_l246_42) begin
          _zz_io_push_payload_wstrb[43 : 40] = 4'b1111;
        end
        if(when_MemoryEngine_l246_43) begin
          _zz_io_push_payload_wstrb[47 : 44] = 4'b1111;
        end
        if(when_MemoryEngine_l246_44) begin
          _zz_io_push_payload_wstrb[51 : 48] = 4'b1111;
        end
        if(when_MemoryEngine_l246_45) begin
          _zz_io_push_payload_wstrb[55 : 52] = 4'b1111;
        end
        if(when_MemoryEngine_l246_46) begin
          _zz_io_push_payload_wstrb[59 : 56] = 4'b1111;
        end
        if(when_MemoryEngine_l246_47) begin
          _zz_io_push_payload_wstrb[63 : 60] = 4'b1111;
        end
        if(when_MemoryEngine_l246_48) begin
          _zz_io_push_payload_wstrb[3 : 0] = 4'b1111;
        end
        if(when_MemoryEngine_l246_49) begin
          _zz_io_push_payload_wstrb[7 : 4] = 4'b1111;
        end
        if(when_MemoryEngine_l246_50) begin
          _zz_io_push_payload_wstrb[11 : 8] = 4'b1111;
        end
        if(when_MemoryEngine_l246_51) begin
          _zz_io_push_payload_wstrb[15 : 12] = 4'b1111;
        end
        if(when_MemoryEngine_l246_52) begin
          _zz_io_push_payload_wstrb[19 : 16] = 4'b1111;
        end
        if(when_MemoryEngine_l246_53) begin
          _zz_io_push_payload_wstrb[23 : 20] = 4'b1111;
        end
        if(when_MemoryEngine_l246_54) begin
          _zz_io_push_payload_wstrb[27 : 24] = 4'b1111;
        end
        if(when_MemoryEngine_l246_55) begin
          _zz_io_push_payload_wstrb[31 : 28] = 4'b1111;
        end
        if(when_MemoryEngine_l246_56) begin
          _zz_io_push_payload_wstrb[35 : 32] = 4'b1111;
        end
        if(when_MemoryEngine_l246_57) begin
          _zz_io_push_payload_wstrb[39 : 36] = 4'b1111;
        end
        if(when_MemoryEngine_l246_58) begin
          _zz_io_push_payload_wstrb[43 : 40] = 4'b1111;
        end
        if(when_MemoryEngine_l246_59) begin
          _zz_io_push_payload_wstrb[47 : 44] = 4'b1111;
        end
        if(when_MemoryEngine_l246_60) begin
          _zz_io_push_payload_wstrb[51 : 48] = 4'b1111;
        end
        if(when_MemoryEngine_l246_61) begin
          _zz_io_push_payload_wstrb[55 : 52] = 4'b1111;
        end
        if(when_MemoryEngine_l246_62) begin
          _zz_io_push_payload_wstrb[59 : 56] = 4'b1111;
        end
        if(when_MemoryEngine_l246_63) begin
          _zz_io_push_payload_wstrb[63 : 60] = 4'b1111;
        end
        if(when_MemoryEngine_l246_64) begin
          _zz_io_push_payload_wstrb[3 : 0] = 4'b1111;
        end
        if(when_MemoryEngine_l246_65) begin
          _zz_io_push_payload_wstrb[7 : 4] = 4'b1111;
        end
        if(when_MemoryEngine_l246_66) begin
          _zz_io_push_payload_wstrb[11 : 8] = 4'b1111;
        end
        if(when_MemoryEngine_l246_67) begin
          _zz_io_push_payload_wstrb[15 : 12] = 4'b1111;
        end
        if(when_MemoryEngine_l246_68) begin
          _zz_io_push_payload_wstrb[19 : 16] = 4'b1111;
        end
        if(when_MemoryEngine_l246_69) begin
          _zz_io_push_payload_wstrb[23 : 20] = 4'b1111;
        end
        if(when_MemoryEngine_l246_70) begin
          _zz_io_push_payload_wstrb[27 : 24] = 4'b1111;
        end
        if(when_MemoryEngine_l246_71) begin
          _zz_io_push_payload_wstrb[31 : 28] = 4'b1111;
        end
        if(when_MemoryEngine_l246_72) begin
          _zz_io_push_payload_wstrb[35 : 32] = 4'b1111;
        end
        if(when_MemoryEngine_l246_73) begin
          _zz_io_push_payload_wstrb[39 : 36] = 4'b1111;
        end
        if(when_MemoryEngine_l246_74) begin
          _zz_io_push_payload_wstrb[43 : 40] = 4'b1111;
        end
        if(when_MemoryEngine_l246_75) begin
          _zz_io_push_payload_wstrb[47 : 44] = 4'b1111;
        end
        if(when_MemoryEngine_l246_76) begin
          _zz_io_push_payload_wstrb[51 : 48] = 4'b1111;
        end
        if(when_MemoryEngine_l246_77) begin
          _zz_io_push_payload_wstrb[55 : 52] = 4'b1111;
        end
        if(when_MemoryEngine_l246_78) begin
          _zz_io_push_payload_wstrb[59 : 56] = 4'b1111;
        end
        if(when_MemoryEngine_l246_79) begin
          _zz_io_push_payload_wstrb[63 : 60] = 4'b1111;
        end
        if(when_MemoryEngine_l246_80) begin
          _zz_io_push_payload_wstrb[3 : 0] = 4'b1111;
        end
        if(when_MemoryEngine_l246_81) begin
          _zz_io_push_payload_wstrb[7 : 4] = 4'b1111;
        end
        if(when_MemoryEngine_l246_82) begin
          _zz_io_push_payload_wstrb[11 : 8] = 4'b1111;
        end
        if(when_MemoryEngine_l246_83) begin
          _zz_io_push_payload_wstrb[15 : 12] = 4'b1111;
        end
        if(when_MemoryEngine_l246_84) begin
          _zz_io_push_payload_wstrb[19 : 16] = 4'b1111;
        end
        if(when_MemoryEngine_l246_85) begin
          _zz_io_push_payload_wstrb[23 : 20] = 4'b1111;
        end
        if(when_MemoryEngine_l246_86) begin
          _zz_io_push_payload_wstrb[27 : 24] = 4'b1111;
        end
        if(when_MemoryEngine_l246_87) begin
          _zz_io_push_payload_wstrb[31 : 28] = 4'b1111;
        end
        if(when_MemoryEngine_l246_88) begin
          _zz_io_push_payload_wstrb[35 : 32] = 4'b1111;
        end
        if(when_MemoryEngine_l246_89) begin
          _zz_io_push_payload_wstrb[39 : 36] = 4'b1111;
        end
        if(when_MemoryEngine_l246_90) begin
          _zz_io_push_payload_wstrb[43 : 40] = 4'b1111;
        end
        if(when_MemoryEngine_l246_91) begin
          _zz_io_push_payload_wstrb[47 : 44] = 4'b1111;
        end
        if(when_MemoryEngine_l246_92) begin
          _zz_io_push_payload_wstrb[51 : 48] = 4'b1111;
        end
        if(when_MemoryEngine_l246_93) begin
          _zz_io_push_payload_wstrb[55 : 52] = 4'b1111;
        end
        if(when_MemoryEngine_l246_94) begin
          _zz_io_push_payload_wstrb[59 : 56] = 4'b1111;
        end
        if(when_MemoryEngine_l246_95) begin
          _zz_io_push_payload_wstrb[63 : 60] = 4'b1111;
        end
        if(when_MemoryEngine_l246_96) begin
          _zz_io_push_payload_wstrb[3 : 0] = 4'b1111;
        end
        if(when_MemoryEngine_l246_97) begin
          _zz_io_push_payload_wstrb[7 : 4] = 4'b1111;
        end
        if(when_MemoryEngine_l246_98) begin
          _zz_io_push_payload_wstrb[11 : 8] = 4'b1111;
        end
        if(when_MemoryEngine_l246_99) begin
          _zz_io_push_payload_wstrb[15 : 12] = 4'b1111;
        end
        if(when_MemoryEngine_l246_100) begin
          _zz_io_push_payload_wstrb[19 : 16] = 4'b1111;
        end
        if(when_MemoryEngine_l246_101) begin
          _zz_io_push_payload_wstrb[23 : 20] = 4'b1111;
        end
        if(when_MemoryEngine_l246_102) begin
          _zz_io_push_payload_wstrb[27 : 24] = 4'b1111;
        end
        if(when_MemoryEngine_l246_103) begin
          _zz_io_push_payload_wstrb[31 : 28] = 4'b1111;
        end
        if(when_MemoryEngine_l246_104) begin
          _zz_io_push_payload_wstrb[35 : 32] = 4'b1111;
        end
        if(when_MemoryEngine_l246_105) begin
          _zz_io_push_payload_wstrb[39 : 36] = 4'b1111;
        end
        if(when_MemoryEngine_l246_106) begin
          _zz_io_push_payload_wstrb[43 : 40] = 4'b1111;
        end
        if(when_MemoryEngine_l246_107) begin
          _zz_io_push_payload_wstrb[47 : 44] = 4'b1111;
        end
        if(when_MemoryEngine_l246_108) begin
          _zz_io_push_payload_wstrb[51 : 48] = 4'b1111;
        end
        if(when_MemoryEngine_l246_109) begin
          _zz_io_push_payload_wstrb[55 : 52] = 4'b1111;
        end
        if(when_MemoryEngine_l246_110) begin
          _zz_io_push_payload_wstrb[59 : 56] = 4'b1111;
        end
        if(when_MemoryEngine_l246_111) begin
          _zz_io_push_payload_wstrb[63 : 60] = 4'b1111;
        end
        if(when_MemoryEngine_l246_112) begin
          _zz_io_push_payload_wstrb[3 : 0] = 4'b1111;
        end
        if(when_MemoryEngine_l246_113) begin
          _zz_io_push_payload_wstrb[7 : 4] = 4'b1111;
        end
        if(when_MemoryEngine_l246_114) begin
          _zz_io_push_payload_wstrb[11 : 8] = 4'b1111;
        end
        if(when_MemoryEngine_l246_115) begin
          _zz_io_push_payload_wstrb[15 : 12] = 4'b1111;
        end
        if(when_MemoryEngine_l246_116) begin
          _zz_io_push_payload_wstrb[19 : 16] = 4'b1111;
        end
        if(when_MemoryEngine_l246_117) begin
          _zz_io_push_payload_wstrb[23 : 20] = 4'b1111;
        end
        if(when_MemoryEngine_l246_118) begin
          _zz_io_push_payload_wstrb[27 : 24] = 4'b1111;
        end
        if(when_MemoryEngine_l246_119) begin
          _zz_io_push_payload_wstrb[31 : 28] = 4'b1111;
        end
        if(when_MemoryEngine_l246_120) begin
          _zz_io_push_payload_wstrb[35 : 32] = 4'b1111;
        end
        if(when_MemoryEngine_l246_121) begin
          _zz_io_push_payload_wstrb[39 : 36] = 4'b1111;
        end
        if(when_MemoryEngine_l246_122) begin
          _zz_io_push_payload_wstrb[43 : 40] = 4'b1111;
        end
        if(when_MemoryEngine_l246_123) begin
          _zz_io_push_payload_wstrb[47 : 44] = 4'b1111;
        end
        if(when_MemoryEngine_l246_124) begin
          _zz_io_push_payload_wstrb[51 : 48] = 4'b1111;
        end
        if(when_MemoryEngine_l246_125) begin
          _zz_io_push_payload_wstrb[55 : 52] = 4'b1111;
        end
        if(when_MemoryEngine_l246_126) begin
          _zz_io_push_payload_wstrb[59 : 56] = 4'b1111;
        end
        if(when_MemoryEngine_l246_127) begin
          _zz_io_push_payload_wstrb[63 : 60] = 4'b1111;
        end
      end
      default : begin
      end
    endcase
  end

  assign when_MemoryEngine_l235 = (_zz_when_MemoryEngine_l235 == 4'b0000);
  assign when_MemoryEngine_l235_1 = (_zz_when_MemoryEngine_l235 == 4'b0001);
  assign when_MemoryEngine_l235_2 = (_zz_when_MemoryEngine_l235 == 4'b0010);
  assign when_MemoryEngine_l235_3 = (_zz_when_MemoryEngine_l235 == 4'b0011);
  assign when_MemoryEngine_l235_4 = (_zz_when_MemoryEngine_l235 == 4'b0100);
  assign when_MemoryEngine_l235_5 = (_zz_when_MemoryEngine_l235 == 4'b0101);
  assign when_MemoryEngine_l235_6 = (_zz_when_MemoryEngine_l235 == 4'b0110);
  assign when_MemoryEngine_l235_7 = (_zz_when_MemoryEngine_l235 == 4'b0111);
  assign when_MemoryEngine_l235_8 = (_zz_when_MemoryEngine_l235 == 4'b1000);
  assign when_MemoryEngine_l235_9 = (_zz_when_MemoryEngine_l235 == 4'b1001);
  assign when_MemoryEngine_l235_10 = (_zz_when_MemoryEngine_l235 == 4'b1010);
  assign when_MemoryEngine_l235_11 = (_zz_when_MemoryEngine_l235 == 4'b1011);
  assign when_MemoryEngine_l235_12 = (_zz_when_MemoryEngine_l235 == 4'b1100);
  assign when_MemoryEngine_l235_13 = (_zz_when_MemoryEngine_l235 == 4'b1101);
  assign when_MemoryEngine_l235_14 = (_zz_when_MemoryEngine_l235 == 4'b1110);
  assign when_MemoryEngine_l235_15 = (_zz_when_MemoryEngine_l235 == 4'b1111);
  assign _zz_when_MemoryEngine_l246 = (_zz_when_MemoryEngine_l235 + 4'b0000);
  assign when_MemoryEngine_l246 = (_zz_when_MemoryEngine_l246 == 4'b0000);
  assign when_MemoryEngine_l246_1 = (_zz_when_MemoryEngine_l246 == 4'b0001);
  assign when_MemoryEngine_l246_2 = (_zz_when_MemoryEngine_l246 == 4'b0010);
  assign when_MemoryEngine_l246_3 = (_zz_when_MemoryEngine_l246 == 4'b0011);
  assign when_MemoryEngine_l246_4 = (_zz_when_MemoryEngine_l246 == 4'b0100);
  assign when_MemoryEngine_l246_5 = (_zz_when_MemoryEngine_l246 == 4'b0101);
  assign when_MemoryEngine_l246_6 = (_zz_when_MemoryEngine_l246 == 4'b0110);
  assign when_MemoryEngine_l246_7 = (_zz_when_MemoryEngine_l246 == 4'b0111);
  assign when_MemoryEngine_l246_8 = (_zz_when_MemoryEngine_l246 == 4'b1000);
  assign when_MemoryEngine_l246_9 = (_zz_when_MemoryEngine_l246 == 4'b1001);
  assign when_MemoryEngine_l246_10 = (_zz_when_MemoryEngine_l246 == 4'b1010);
  assign when_MemoryEngine_l246_11 = (_zz_when_MemoryEngine_l246 == 4'b1011);
  assign when_MemoryEngine_l246_12 = (_zz_when_MemoryEngine_l246 == 4'b1100);
  assign when_MemoryEngine_l246_13 = (_zz_when_MemoryEngine_l246 == 4'b1101);
  assign when_MemoryEngine_l246_14 = (_zz_when_MemoryEngine_l246 == 4'b1110);
  assign when_MemoryEngine_l246_15 = (_zz_when_MemoryEngine_l246 == 4'b1111);
  assign _zz_when_MemoryEngine_l246_1 = (_zz_when_MemoryEngine_l235 + 4'b0001);
  assign when_MemoryEngine_l246_16 = (_zz_when_MemoryEngine_l246_1 == 4'b0000);
  assign when_MemoryEngine_l246_17 = (_zz_when_MemoryEngine_l246_1 == 4'b0001);
  assign when_MemoryEngine_l246_18 = (_zz_when_MemoryEngine_l246_1 == 4'b0010);
  assign when_MemoryEngine_l246_19 = (_zz_when_MemoryEngine_l246_1 == 4'b0011);
  assign when_MemoryEngine_l246_20 = (_zz_when_MemoryEngine_l246_1 == 4'b0100);
  assign when_MemoryEngine_l246_21 = (_zz_when_MemoryEngine_l246_1 == 4'b0101);
  assign when_MemoryEngine_l246_22 = (_zz_when_MemoryEngine_l246_1 == 4'b0110);
  assign when_MemoryEngine_l246_23 = (_zz_when_MemoryEngine_l246_1 == 4'b0111);
  assign when_MemoryEngine_l246_24 = (_zz_when_MemoryEngine_l246_1 == 4'b1000);
  assign when_MemoryEngine_l246_25 = (_zz_when_MemoryEngine_l246_1 == 4'b1001);
  assign when_MemoryEngine_l246_26 = (_zz_when_MemoryEngine_l246_1 == 4'b1010);
  assign when_MemoryEngine_l246_27 = (_zz_when_MemoryEngine_l246_1 == 4'b1011);
  assign when_MemoryEngine_l246_28 = (_zz_when_MemoryEngine_l246_1 == 4'b1100);
  assign when_MemoryEngine_l246_29 = (_zz_when_MemoryEngine_l246_1 == 4'b1101);
  assign when_MemoryEngine_l246_30 = (_zz_when_MemoryEngine_l246_1 == 4'b1110);
  assign when_MemoryEngine_l246_31 = (_zz_when_MemoryEngine_l246_1 == 4'b1111);
  assign _zz_when_MemoryEngine_l246_2 = (_zz_when_MemoryEngine_l235 + 4'b0010);
  assign when_MemoryEngine_l246_32 = (_zz_when_MemoryEngine_l246_2 == 4'b0000);
  assign when_MemoryEngine_l246_33 = (_zz_when_MemoryEngine_l246_2 == 4'b0001);
  assign when_MemoryEngine_l246_34 = (_zz_when_MemoryEngine_l246_2 == 4'b0010);
  assign when_MemoryEngine_l246_35 = (_zz_when_MemoryEngine_l246_2 == 4'b0011);
  assign when_MemoryEngine_l246_36 = (_zz_when_MemoryEngine_l246_2 == 4'b0100);
  assign when_MemoryEngine_l246_37 = (_zz_when_MemoryEngine_l246_2 == 4'b0101);
  assign when_MemoryEngine_l246_38 = (_zz_when_MemoryEngine_l246_2 == 4'b0110);
  assign when_MemoryEngine_l246_39 = (_zz_when_MemoryEngine_l246_2 == 4'b0111);
  assign when_MemoryEngine_l246_40 = (_zz_when_MemoryEngine_l246_2 == 4'b1000);
  assign when_MemoryEngine_l246_41 = (_zz_when_MemoryEngine_l246_2 == 4'b1001);
  assign when_MemoryEngine_l246_42 = (_zz_when_MemoryEngine_l246_2 == 4'b1010);
  assign when_MemoryEngine_l246_43 = (_zz_when_MemoryEngine_l246_2 == 4'b1011);
  assign when_MemoryEngine_l246_44 = (_zz_when_MemoryEngine_l246_2 == 4'b1100);
  assign when_MemoryEngine_l246_45 = (_zz_when_MemoryEngine_l246_2 == 4'b1101);
  assign when_MemoryEngine_l246_46 = (_zz_when_MemoryEngine_l246_2 == 4'b1110);
  assign when_MemoryEngine_l246_47 = (_zz_when_MemoryEngine_l246_2 == 4'b1111);
  assign _zz_when_MemoryEngine_l246_3 = (_zz_when_MemoryEngine_l235 + 4'b0011);
  assign when_MemoryEngine_l246_48 = (_zz_when_MemoryEngine_l246_3 == 4'b0000);
  assign when_MemoryEngine_l246_49 = (_zz_when_MemoryEngine_l246_3 == 4'b0001);
  assign when_MemoryEngine_l246_50 = (_zz_when_MemoryEngine_l246_3 == 4'b0010);
  assign when_MemoryEngine_l246_51 = (_zz_when_MemoryEngine_l246_3 == 4'b0011);
  assign when_MemoryEngine_l246_52 = (_zz_when_MemoryEngine_l246_3 == 4'b0100);
  assign when_MemoryEngine_l246_53 = (_zz_when_MemoryEngine_l246_3 == 4'b0101);
  assign when_MemoryEngine_l246_54 = (_zz_when_MemoryEngine_l246_3 == 4'b0110);
  assign when_MemoryEngine_l246_55 = (_zz_when_MemoryEngine_l246_3 == 4'b0111);
  assign when_MemoryEngine_l246_56 = (_zz_when_MemoryEngine_l246_3 == 4'b1000);
  assign when_MemoryEngine_l246_57 = (_zz_when_MemoryEngine_l246_3 == 4'b1001);
  assign when_MemoryEngine_l246_58 = (_zz_when_MemoryEngine_l246_3 == 4'b1010);
  assign when_MemoryEngine_l246_59 = (_zz_when_MemoryEngine_l246_3 == 4'b1011);
  assign when_MemoryEngine_l246_60 = (_zz_when_MemoryEngine_l246_3 == 4'b1100);
  assign when_MemoryEngine_l246_61 = (_zz_when_MemoryEngine_l246_3 == 4'b1101);
  assign when_MemoryEngine_l246_62 = (_zz_when_MemoryEngine_l246_3 == 4'b1110);
  assign when_MemoryEngine_l246_63 = (_zz_when_MemoryEngine_l246_3 == 4'b1111);
  assign _zz_when_MemoryEngine_l246_4 = (_zz_when_MemoryEngine_l235 + 4'b0100);
  assign when_MemoryEngine_l246_64 = (_zz_when_MemoryEngine_l246_4 == 4'b0000);
  assign when_MemoryEngine_l246_65 = (_zz_when_MemoryEngine_l246_4 == 4'b0001);
  assign when_MemoryEngine_l246_66 = (_zz_when_MemoryEngine_l246_4 == 4'b0010);
  assign when_MemoryEngine_l246_67 = (_zz_when_MemoryEngine_l246_4 == 4'b0011);
  assign when_MemoryEngine_l246_68 = (_zz_when_MemoryEngine_l246_4 == 4'b0100);
  assign when_MemoryEngine_l246_69 = (_zz_when_MemoryEngine_l246_4 == 4'b0101);
  assign when_MemoryEngine_l246_70 = (_zz_when_MemoryEngine_l246_4 == 4'b0110);
  assign when_MemoryEngine_l246_71 = (_zz_when_MemoryEngine_l246_4 == 4'b0111);
  assign when_MemoryEngine_l246_72 = (_zz_when_MemoryEngine_l246_4 == 4'b1000);
  assign when_MemoryEngine_l246_73 = (_zz_when_MemoryEngine_l246_4 == 4'b1001);
  assign when_MemoryEngine_l246_74 = (_zz_when_MemoryEngine_l246_4 == 4'b1010);
  assign when_MemoryEngine_l246_75 = (_zz_when_MemoryEngine_l246_4 == 4'b1011);
  assign when_MemoryEngine_l246_76 = (_zz_when_MemoryEngine_l246_4 == 4'b1100);
  assign when_MemoryEngine_l246_77 = (_zz_when_MemoryEngine_l246_4 == 4'b1101);
  assign when_MemoryEngine_l246_78 = (_zz_when_MemoryEngine_l246_4 == 4'b1110);
  assign when_MemoryEngine_l246_79 = (_zz_when_MemoryEngine_l246_4 == 4'b1111);
  assign _zz_when_MemoryEngine_l246_5 = (_zz_when_MemoryEngine_l235 + 4'b0101);
  assign when_MemoryEngine_l246_80 = (_zz_when_MemoryEngine_l246_5 == 4'b0000);
  assign when_MemoryEngine_l246_81 = (_zz_when_MemoryEngine_l246_5 == 4'b0001);
  assign when_MemoryEngine_l246_82 = (_zz_when_MemoryEngine_l246_5 == 4'b0010);
  assign when_MemoryEngine_l246_83 = (_zz_when_MemoryEngine_l246_5 == 4'b0011);
  assign when_MemoryEngine_l246_84 = (_zz_when_MemoryEngine_l246_5 == 4'b0100);
  assign when_MemoryEngine_l246_85 = (_zz_when_MemoryEngine_l246_5 == 4'b0101);
  assign when_MemoryEngine_l246_86 = (_zz_when_MemoryEngine_l246_5 == 4'b0110);
  assign when_MemoryEngine_l246_87 = (_zz_when_MemoryEngine_l246_5 == 4'b0111);
  assign when_MemoryEngine_l246_88 = (_zz_when_MemoryEngine_l246_5 == 4'b1000);
  assign when_MemoryEngine_l246_89 = (_zz_when_MemoryEngine_l246_5 == 4'b1001);
  assign when_MemoryEngine_l246_90 = (_zz_when_MemoryEngine_l246_5 == 4'b1010);
  assign when_MemoryEngine_l246_91 = (_zz_when_MemoryEngine_l246_5 == 4'b1011);
  assign when_MemoryEngine_l246_92 = (_zz_when_MemoryEngine_l246_5 == 4'b1100);
  assign when_MemoryEngine_l246_93 = (_zz_when_MemoryEngine_l246_5 == 4'b1101);
  assign when_MemoryEngine_l246_94 = (_zz_when_MemoryEngine_l246_5 == 4'b1110);
  assign when_MemoryEngine_l246_95 = (_zz_when_MemoryEngine_l246_5 == 4'b1111);
  assign _zz_when_MemoryEngine_l246_6 = (_zz_when_MemoryEngine_l235 + 4'b0110);
  assign when_MemoryEngine_l246_96 = (_zz_when_MemoryEngine_l246_6 == 4'b0000);
  assign when_MemoryEngine_l246_97 = (_zz_when_MemoryEngine_l246_6 == 4'b0001);
  assign when_MemoryEngine_l246_98 = (_zz_when_MemoryEngine_l246_6 == 4'b0010);
  assign when_MemoryEngine_l246_99 = (_zz_when_MemoryEngine_l246_6 == 4'b0011);
  assign when_MemoryEngine_l246_100 = (_zz_when_MemoryEngine_l246_6 == 4'b0100);
  assign when_MemoryEngine_l246_101 = (_zz_when_MemoryEngine_l246_6 == 4'b0101);
  assign when_MemoryEngine_l246_102 = (_zz_when_MemoryEngine_l246_6 == 4'b0110);
  assign when_MemoryEngine_l246_103 = (_zz_when_MemoryEngine_l246_6 == 4'b0111);
  assign when_MemoryEngine_l246_104 = (_zz_when_MemoryEngine_l246_6 == 4'b1000);
  assign when_MemoryEngine_l246_105 = (_zz_when_MemoryEngine_l246_6 == 4'b1001);
  assign when_MemoryEngine_l246_106 = (_zz_when_MemoryEngine_l246_6 == 4'b1010);
  assign when_MemoryEngine_l246_107 = (_zz_when_MemoryEngine_l246_6 == 4'b1011);
  assign when_MemoryEngine_l246_108 = (_zz_when_MemoryEngine_l246_6 == 4'b1100);
  assign when_MemoryEngine_l246_109 = (_zz_when_MemoryEngine_l246_6 == 4'b1101);
  assign when_MemoryEngine_l246_110 = (_zz_when_MemoryEngine_l246_6 == 4'b1110);
  assign when_MemoryEngine_l246_111 = (_zz_when_MemoryEngine_l246_6 == 4'b1111);
  assign _zz_when_MemoryEngine_l246_7 = (_zz_when_MemoryEngine_l235 + 4'b0111);
  assign when_MemoryEngine_l246_112 = (_zz_when_MemoryEngine_l246_7 == 4'b0000);
  assign when_MemoryEngine_l246_113 = (_zz_when_MemoryEngine_l246_7 == 4'b0001);
  assign when_MemoryEngine_l246_114 = (_zz_when_MemoryEngine_l246_7 == 4'b0010);
  assign when_MemoryEngine_l246_115 = (_zz_when_MemoryEngine_l246_7 == 4'b0011);
  assign when_MemoryEngine_l246_116 = (_zz_when_MemoryEngine_l246_7 == 4'b0100);
  assign when_MemoryEngine_l246_117 = (_zz_when_MemoryEngine_l246_7 == 4'b0101);
  assign when_MemoryEngine_l246_118 = (_zz_when_MemoryEngine_l246_7 == 4'b0110);
  assign when_MemoryEngine_l246_119 = (_zz_when_MemoryEngine_l246_7 == 4'b0111);
  assign when_MemoryEngine_l246_120 = (_zz_when_MemoryEngine_l246_7 == 4'b1000);
  assign when_MemoryEngine_l246_121 = (_zz_when_MemoryEngine_l246_7 == 4'b1001);
  assign when_MemoryEngine_l246_122 = (_zz_when_MemoryEngine_l246_7 == 4'b1010);
  assign when_MemoryEngine_l246_123 = (_zz_when_MemoryEngine_l246_7 == 4'b1011);
  assign when_MemoryEngine_l246_124 = (_zz_when_MemoryEngine_l246_7 == 4'b1100);
  assign when_MemoryEngine_l246_125 = (_zz_when_MemoryEngine_l246_7 == 4'b1101);
  assign when_MemoryEngine_l246_126 = (_zz_when_MemoryEngine_l246_7 == 4'b1110);
  assign when_MemoryEngine_l246_127 = (_zz_when_MemoryEngine_l246_7 == 4'b1111);
  always @(*) begin
    storeReqFifo_io_pop_ready = 1'b0;
    case(state)
      MemState_IDLE : begin
        if(storeReqFifo_io_pop_valid) begin
          storeReqFifo_io_pop_ready = 1'b1;
        end
      end
      MemState_STORE_AW_W : begin
      end
      default : begin
      end
    endcase
  end

  assign io_axiMaster_ar_valid = loadReqValid;
  assign io_axiMaster_ar_payload_addr = loadReqEntry_axiAddr;
  assign io_axiMaster_ar_payload_len = 8'h0;
  assign io_axiMaster_ar_payload_size = axiSizeVal;
  assign io_axiMaster_ar_payload_burst = 2'b01;
  assign io_axiMaster_ar_payload_id = 4'b0000;
  assign io_axiMaster_r_ready = loadReqValid;
  assign when_MemoryEngine_l285 = (io_axiMaster_r_valid && loadReqValid);
  assign when_MemoryEngine_l291 = (loadReqEntry_slotIdx == 1'b0);
  assign when_MemoryEngine_l292 = (! loadReqEntry_isVector);
  always @(*) begin
    _zz_io_loadWriteReqs_0_payload_data = 32'h0;
    if(when_MemoryEngine_l297) begin
      _zz_io_loadWriteReqs_0_payload_data = io_axiMaster_r_payload_data[31 : 0];
    end
    if(when_MemoryEngine_l297_1) begin
      _zz_io_loadWriteReqs_0_payload_data = io_axiMaster_r_payload_data[63 : 32];
    end
    if(when_MemoryEngine_l297_2) begin
      _zz_io_loadWriteReqs_0_payload_data = io_axiMaster_r_payload_data[95 : 64];
    end
    if(when_MemoryEngine_l297_3) begin
      _zz_io_loadWriteReqs_0_payload_data = io_axiMaster_r_payload_data[127 : 96];
    end
    if(when_MemoryEngine_l297_4) begin
      _zz_io_loadWriteReqs_0_payload_data = io_axiMaster_r_payload_data[159 : 128];
    end
    if(when_MemoryEngine_l297_5) begin
      _zz_io_loadWriteReqs_0_payload_data = io_axiMaster_r_payload_data[191 : 160];
    end
    if(when_MemoryEngine_l297_6) begin
      _zz_io_loadWriteReqs_0_payload_data = io_axiMaster_r_payload_data[223 : 192];
    end
    if(when_MemoryEngine_l297_7) begin
      _zz_io_loadWriteReqs_0_payload_data = io_axiMaster_r_payload_data[255 : 224];
    end
    if(when_MemoryEngine_l297_8) begin
      _zz_io_loadWriteReqs_0_payload_data = io_axiMaster_r_payload_data[287 : 256];
    end
    if(when_MemoryEngine_l297_9) begin
      _zz_io_loadWriteReqs_0_payload_data = io_axiMaster_r_payload_data[319 : 288];
    end
    if(when_MemoryEngine_l297_10) begin
      _zz_io_loadWriteReqs_0_payload_data = io_axiMaster_r_payload_data[351 : 320];
    end
    if(when_MemoryEngine_l297_11) begin
      _zz_io_loadWriteReqs_0_payload_data = io_axiMaster_r_payload_data[383 : 352];
    end
    if(when_MemoryEngine_l297_12) begin
      _zz_io_loadWriteReqs_0_payload_data = io_axiMaster_r_payload_data[415 : 384];
    end
    if(when_MemoryEngine_l297_13) begin
      _zz_io_loadWriteReqs_0_payload_data = io_axiMaster_r_payload_data[447 : 416];
    end
    if(when_MemoryEngine_l297_14) begin
      _zz_io_loadWriteReqs_0_payload_data = io_axiMaster_r_payload_data[479 : 448];
    end
    if(when_MemoryEngine_l297_15) begin
      _zz_io_loadWriteReqs_0_payload_data = io_axiMaster_r_payload_data[511 : 480];
    end
  end

  assign when_MemoryEngine_l297 = (loadReqEntry_wordOff == 4'b0000);
  assign when_MemoryEngine_l297_1 = (loadReqEntry_wordOff == 4'b0001);
  assign when_MemoryEngine_l297_2 = (loadReqEntry_wordOff == 4'b0010);
  assign when_MemoryEngine_l297_3 = (loadReqEntry_wordOff == 4'b0011);
  assign when_MemoryEngine_l297_4 = (loadReqEntry_wordOff == 4'b0100);
  assign when_MemoryEngine_l297_5 = (loadReqEntry_wordOff == 4'b0101);
  assign when_MemoryEngine_l297_6 = (loadReqEntry_wordOff == 4'b0110);
  assign when_MemoryEngine_l297_7 = (loadReqEntry_wordOff == 4'b0111);
  assign when_MemoryEngine_l297_8 = (loadReqEntry_wordOff == 4'b1000);
  assign when_MemoryEngine_l297_9 = (loadReqEntry_wordOff == 4'b1001);
  assign when_MemoryEngine_l297_10 = (loadReqEntry_wordOff == 4'b1010);
  assign when_MemoryEngine_l297_11 = (loadReqEntry_wordOff == 4'b1011);
  assign when_MemoryEngine_l297_12 = (loadReqEntry_wordOff == 4'b1100);
  assign when_MemoryEngine_l297_13 = (loadReqEntry_wordOff == 4'b1101);
  assign when_MemoryEngine_l297_14 = (loadReqEntry_wordOff == 4'b1110);
  assign when_MemoryEngine_l297_15 = (loadReqEntry_wordOff == 4'b1111);
  always @(*) begin
    _zz_io_vloadWriteReqs_0_0_payload_data = 32'h0;
    if(when_MemoryEngine_l311) begin
      _zz_io_vloadWriteReqs_0_0_payload_data = io_axiMaster_r_payload_data[31 : 0];
    end
    if(when_MemoryEngine_l311_1) begin
      _zz_io_vloadWriteReqs_0_0_payload_data = io_axiMaster_r_payload_data[63 : 32];
    end
    if(when_MemoryEngine_l311_2) begin
      _zz_io_vloadWriteReqs_0_0_payload_data = io_axiMaster_r_payload_data[95 : 64];
    end
    if(when_MemoryEngine_l311_3) begin
      _zz_io_vloadWriteReqs_0_0_payload_data = io_axiMaster_r_payload_data[127 : 96];
    end
    if(when_MemoryEngine_l311_4) begin
      _zz_io_vloadWriteReqs_0_0_payload_data = io_axiMaster_r_payload_data[159 : 128];
    end
    if(when_MemoryEngine_l311_5) begin
      _zz_io_vloadWriteReqs_0_0_payload_data = io_axiMaster_r_payload_data[191 : 160];
    end
    if(when_MemoryEngine_l311_6) begin
      _zz_io_vloadWriteReqs_0_0_payload_data = io_axiMaster_r_payload_data[223 : 192];
    end
    if(when_MemoryEngine_l311_7) begin
      _zz_io_vloadWriteReqs_0_0_payload_data = io_axiMaster_r_payload_data[255 : 224];
    end
    if(when_MemoryEngine_l311_8) begin
      _zz_io_vloadWriteReqs_0_0_payload_data = io_axiMaster_r_payload_data[287 : 256];
    end
    if(when_MemoryEngine_l311_9) begin
      _zz_io_vloadWriteReqs_0_0_payload_data = io_axiMaster_r_payload_data[319 : 288];
    end
    if(when_MemoryEngine_l311_10) begin
      _zz_io_vloadWriteReqs_0_0_payload_data = io_axiMaster_r_payload_data[351 : 320];
    end
    if(when_MemoryEngine_l311_11) begin
      _zz_io_vloadWriteReqs_0_0_payload_data = io_axiMaster_r_payload_data[383 : 352];
    end
    if(when_MemoryEngine_l311_12) begin
      _zz_io_vloadWriteReqs_0_0_payload_data = io_axiMaster_r_payload_data[415 : 384];
    end
    if(when_MemoryEngine_l311_13) begin
      _zz_io_vloadWriteReqs_0_0_payload_data = io_axiMaster_r_payload_data[447 : 416];
    end
    if(when_MemoryEngine_l311_14) begin
      _zz_io_vloadWriteReqs_0_0_payload_data = io_axiMaster_r_payload_data[479 : 448];
    end
    if(when_MemoryEngine_l311_15) begin
      _zz_io_vloadWriteReqs_0_0_payload_data = io_axiMaster_r_payload_data[511 : 480];
    end
  end

  assign _zz_when_MemoryEngine_l311 = (loadReqEntry_wordOff + 4'b0000);
  assign when_MemoryEngine_l311 = (_zz_when_MemoryEngine_l311 == 4'b0000);
  assign when_MemoryEngine_l311_1 = (_zz_when_MemoryEngine_l311 == 4'b0001);
  assign when_MemoryEngine_l311_2 = (_zz_when_MemoryEngine_l311 == 4'b0010);
  assign when_MemoryEngine_l311_3 = (_zz_when_MemoryEngine_l311 == 4'b0011);
  assign when_MemoryEngine_l311_4 = (_zz_when_MemoryEngine_l311 == 4'b0100);
  assign when_MemoryEngine_l311_5 = (_zz_when_MemoryEngine_l311 == 4'b0101);
  assign when_MemoryEngine_l311_6 = (_zz_when_MemoryEngine_l311 == 4'b0110);
  assign when_MemoryEngine_l311_7 = (_zz_when_MemoryEngine_l311 == 4'b0111);
  assign when_MemoryEngine_l311_8 = (_zz_when_MemoryEngine_l311 == 4'b1000);
  assign when_MemoryEngine_l311_9 = (_zz_when_MemoryEngine_l311 == 4'b1001);
  assign when_MemoryEngine_l311_10 = (_zz_when_MemoryEngine_l311 == 4'b1010);
  assign when_MemoryEngine_l311_11 = (_zz_when_MemoryEngine_l311 == 4'b1011);
  assign when_MemoryEngine_l311_12 = (_zz_when_MemoryEngine_l311 == 4'b1100);
  assign when_MemoryEngine_l311_13 = (_zz_when_MemoryEngine_l311 == 4'b1101);
  assign when_MemoryEngine_l311_14 = (_zz_when_MemoryEngine_l311 == 4'b1110);
  assign when_MemoryEngine_l311_15 = (_zz_when_MemoryEngine_l311 == 4'b1111);
  always @(*) begin
    _zz_io_vloadWriteReqs_0_1_payload_data = 32'h0;
    if(when_MemoryEngine_l311_16) begin
      _zz_io_vloadWriteReqs_0_1_payload_data = io_axiMaster_r_payload_data[31 : 0];
    end
    if(when_MemoryEngine_l311_17) begin
      _zz_io_vloadWriteReqs_0_1_payload_data = io_axiMaster_r_payload_data[63 : 32];
    end
    if(when_MemoryEngine_l311_18) begin
      _zz_io_vloadWriteReqs_0_1_payload_data = io_axiMaster_r_payload_data[95 : 64];
    end
    if(when_MemoryEngine_l311_19) begin
      _zz_io_vloadWriteReqs_0_1_payload_data = io_axiMaster_r_payload_data[127 : 96];
    end
    if(when_MemoryEngine_l311_20) begin
      _zz_io_vloadWriteReqs_0_1_payload_data = io_axiMaster_r_payload_data[159 : 128];
    end
    if(when_MemoryEngine_l311_21) begin
      _zz_io_vloadWriteReqs_0_1_payload_data = io_axiMaster_r_payload_data[191 : 160];
    end
    if(when_MemoryEngine_l311_22) begin
      _zz_io_vloadWriteReqs_0_1_payload_data = io_axiMaster_r_payload_data[223 : 192];
    end
    if(when_MemoryEngine_l311_23) begin
      _zz_io_vloadWriteReqs_0_1_payload_data = io_axiMaster_r_payload_data[255 : 224];
    end
    if(when_MemoryEngine_l311_24) begin
      _zz_io_vloadWriteReqs_0_1_payload_data = io_axiMaster_r_payload_data[287 : 256];
    end
    if(when_MemoryEngine_l311_25) begin
      _zz_io_vloadWriteReqs_0_1_payload_data = io_axiMaster_r_payload_data[319 : 288];
    end
    if(when_MemoryEngine_l311_26) begin
      _zz_io_vloadWriteReqs_0_1_payload_data = io_axiMaster_r_payload_data[351 : 320];
    end
    if(when_MemoryEngine_l311_27) begin
      _zz_io_vloadWriteReqs_0_1_payload_data = io_axiMaster_r_payload_data[383 : 352];
    end
    if(when_MemoryEngine_l311_28) begin
      _zz_io_vloadWriteReqs_0_1_payload_data = io_axiMaster_r_payload_data[415 : 384];
    end
    if(when_MemoryEngine_l311_29) begin
      _zz_io_vloadWriteReqs_0_1_payload_data = io_axiMaster_r_payload_data[447 : 416];
    end
    if(when_MemoryEngine_l311_30) begin
      _zz_io_vloadWriteReqs_0_1_payload_data = io_axiMaster_r_payload_data[479 : 448];
    end
    if(when_MemoryEngine_l311_31) begin
      _zz_io_vloadWriteReqs_0_1_payload_data = io_axiMaster_r_payload_data[511 : 480];
    end
  end

  assign _zz_when_MemoryEngine_l311_1 = (loadReqEntry_wordOff + 4'b0001);
  assign when_MemoryEngine_l311_16 = (_zz_when_MemoryEngine_l311_1 == 4'b0000);
  assign when_MemoryEngine_l311_17 = (_zz_when_MemoryEngine_l311_1 == 4'b0001);
  assign when_MemoryEngine_l311_18 = (_zz_when_MemoryEngine_l311_1 == 4'b0010);
  assign when_MemoryEngine_l311_19 = (_zz_when_MemoryEngine_l311_1 == 4'b0011);
  assign when_MemoryEngine_l311_20 = (_zz_when_MemoryEngine_l311_1 == 4'b0100);
  assign when_MemoryEngine_l311_21 = (_zz_when_MemoryEngine_l311_1 == 4'b0101);
  assign when_MemoryEngine_l311_22 = (_zz_when_MemoryEngine_l311_1 == 4'b0110);
  assign when_MemoryEngine_l311_23 = (_zz_when_MemoryEngine_l311_1 == 4'b0111);
  assign when_MemoryEngine_l311_24 = (_zz_when_MemoryEngine_l311_1 == 4'b1000);
  assign when_MemoryEngine_l311_25 = (_zz_when_MemoryEngine_l311_1 == 4'b1001);
  assign when_MemoryEngine_l311_26 = (_zz_when_MemoryEngine_l311_1 == 4'b1010);
  assign when_MemoryEngine_l311_27 = (_zz_when_MemoryEngine_l311_1 == 4'b1011);
  assign when_MemoryEngine_l311_28 = (_zz_when_MemoryEngine_l311_1 == 4'b1100);
  assign when_MemoryEngine_l311_29 = (_zz_when_MemoryEngine_l311_1 == 4'b1101);
  assign when_MemoryEngine_l311_30 = (_zz_when_MemoryEngine_l311_1 == 4'b1110);
  assign when_MemoryEngine_l311_31 = (_zz_when_MemoryEngine_l311_1 == 4'b1111);
  always @(*) begin
    _zz_io_vloadWriteReqs_0_2_payload_data = 32'h0;
    if(when_MemoryEngine_l311_32) begin
      _zz_io_vloadWriteReqs_0_2_payload_data = io_axiMaster_r_payload_data[31 : 0];
    end
    if(when_MemoryEngine_l311_33) begin
      _zz_io_vloadWriteReqs_0_2_payload_data = io_axiMaster_r_payload_data[63 : 32];
    end
    if(when_MemoryEngine_l311_34) begin
      _zz_io_vloadWriteReqs_0_2_payload_data = io_axiMaster_r_payload_data[95 : 64];
    end
    if(when_MemoryEngine_l311_35) begin
      _zz_io_vloadWriteReqs_0_2_payload_data = io_axiMaster_r_payload_data[127 : 96];
    end
    if(when_MemoryEngine_l311_36) begin
      _zz_io_vloadWriteReqs_0_2_payload_data = io_axiMaster_r_payload_data[159 : 128];
    end
    if(when_MemoryEngine_l311_37) begin
      _zz_io_vloadWriteReqs_0_2_payload_data = io_axiMaster_r_payload_data[191 : 160];
    end
    if(when_MemoryEngine_l311_38) begin
      _zz_io_vloadWriteReqs_0_2_payload_data = io_axiMaster_r_payload_data[223 : 192];
    end
    if(when_MemoryEngine_l311_39) begin
      _zz_io_vloadWriteReqs_0_2_payload_data = io_axiMaster_r_payload_data[255 : 224];
    end
    if(when_MemoryEngine_l311_40) begin
      _zz_io_vloadWriteReqs_0_2_payload_data = io_axiMaster_r_payload_data[287 : 256];
    end
    if(when_MemoryEngine_l311_41) begin
      _zz_io_vloadWriteReqs_0_2_payload_data = io_axiMaster_r_payload_data[319 : 288];
    end
    if(when_MemoryEngine_l311_42) begin
      _zz_io_vloadWriteReqs_0_2_payload_data = io_axiMaster_r_payload_data[351 : 320];
    end
    if(when_MemoryEngine_l311_43) begin
      _zz_io_vloadWriteReqs_0_2_payload_data = io_axiMaster_r_payload_data[383 : 352];
    end
    if(when_MemoryEngine_l311_44) begin
      _zz_io_vloadWriteReqs_0_2_payload_data = io_axiMaster_r_payload_data[415 : 384];
    end
    if(when_MemoryEngine_l311_45) begin
      _zz_io_vloadWriteReqs_0_2_payload_data = io_axiMaster_r_payload_data[447 : 416];
    end
    if(when_MemoryEngine_l311_46) begin
      _zz_io_vloadWriteReqs_0_2_payload_data = io_axiMaster_r_payload_data[479 : 448];
    end
    if(when_MemoryEngine_l311_47) begin
      _zz_io_vloadWriteReqs_0_2_payload_data = io_axiMaster_r_payload_data[511 : 480];
    end
  end

  assign _zz_when_MemoryEngine_l311_2 = (loadReqEntry_wordOff + 4'b0010);
  assign when_MemoryEngine_l311_32 = (_zz_when_MemoryEngine_l311_2 == 4'b0000);
  assign when_MemoryEngine_l311_33 = (_zz_when_MemoryEngine_l311_2 == 4'b0001);
  assign when_MemoryEngine_l311_34 = (_zz_when_MemoryEngine_l311_2 == 4'b0010);
  assign when_MemoryEngine_l311_35 = (_zz_when_MemoryEngine_l311_2 == 4'b0011);
  assign when_MemoryEngine_l311_36 = (_zz_when_MemoryEngine_l311_2 == 4'b0100);
  assign when_MemoryEngine_l311_37 = (_zz_when_MemoryEngine_l311_2 == 4'b0101);
  assign when_MemoryEngine_l311_38 = (_zz_when_MemoryEngine_l311_2 == 4'b0110);
  assign when_MemoryEngine_l311_39 = (_zz_when_MemoryEngine_l311_2 == 4'b0111);
  assign when_MemoryEngine_l311_40 = (_zz_when_MemoryEngine_l311_2 == 4'b1000);
  assign when_MemoryEngine_l311_41 = (_zz_when_MemoryEngine_l311_2 == 4'b1001);
  assign when_MemoryEngine_l311_42 = (_zz_when_MemoryEngine_l311_2 == 4'b1010);
  assign when_MemoryEngine_l311_43 = (_zz_when_MemoryEngine_l311_2 == 4'b1011);
  assign when_MemoryEngine_l311_44 = (_zz_when_MemoryEngine_l311_2 == 4'b1100);
  assign when_MemoryEngine_l311_45 = (_zz_when_MemoryEngine_l311_2 == 4'b1101);
  assign when_MemoryEngine_l311_46 = (_zz_when_MemoryEngine_l311_2 == 4'b1110);
  assign when_MemoryEngine_l311_47 = (_zz_when_MemoryEngine_l311_2 == 4'b1111);
  always @(*) begin
    _zz_io_vloadWriteReqs_0_3_payload_data = 32'h0;
    if(when_MemoryEngine_l311_48) begin
      _zz_io_vloadWriteReqs_0_3_payload_data = io_axiMaster_r_payload_data[31 : 0];
    end
    if(when_MemoryEngine_l311_49) begin
      _zz_io_vloadWriteReqs_0_3_payload_data = io_axiMaster_r_payload_data[63 : 32];
    end
    if(when_MemoryEngine_l311_50) begin
      _zz_io_vloadWriteReqs_0_3_payload_data = io_axiMaster_r_payload_data[95 : 64];
    end
    if(when_MemoryEngine_l311_51) begin
      _zz_io_vloadWriteReqs_0_3_payload_data = io_axiMaster_r_payload_data[127 : 96];
    end
    if(when_MemoryEngine_l311_52) begin
      _zz_io_vloadWriteReqs_0_3_payload_data = io_axiMaster_r_payload_data[159 : 128];
    end
    if(when_MemoryEngine_l311_53) begin
      _zz_io_vloadWriteReqs_0_3_payload_data = io_axiMaster_r_payload_data[191 : 160];
    end
    if(when_MemoryEngine_l311_54) begin
      _zz_io_vloadWriteReqs_0_3_payload_data = io_axiMaster_r_payload_data[223 : 192];
    end
    if(when_MemoryEngine_l311_55) begin
      _zz_io_vloadWriteReqs_0_3_payload_data = io_axiMaster_r_payload_data[255 : 224];
    end
    if(when_MemoryEngine_l311_56) begin
      _zz_io_vloadWriteReqs_0_3_payload_data = io_axiMaster_r_payload_data[287 : 256];
    end
    if(when_MemoryEngine_l311_57) begin
      _zz_io_vloadWriteReqs_0_3_payload_data = io_axiMaster_r_payload_data[319 : 288];
    end
    if(when_MemoryEngine_l311_58) begin
      _zz_io_vloadWriteReqs_0_3_payload_data = io_axiMaster_r_payload_data[351 : 320];
    end
    if(when_MemoryEngine_l311_59) begin
      _zz_io_vloadWriteReqs_0_3_payload_data = io_axiMaster_r_payload_data[383 : 352];
    end
    if(when_MemoryEngine_l311_60) begin
      _zz_io_vloadWriteReqs_0_3_payload_data = io_axiMaster_r_payload_data[415 : 384];
    end
    if(when_MemoryEngine_l311_61) begin
      _zz_io_vloadWriteReqs_0_3_payload_data = io_axiMaster_r_payload_data[447 : 416];
    end
    if(when_MemoryEngine_l311_62) begin
      _zz_io_vloadWriteReqs_0_3_payload_data = io_axiMaster_r_payload_data[479 : 448];
    end
    if(when_MemoryEngine_l311_63) begin
      _zz_io_vloadWriteReqs_0_3_payload_data = io_axiMaster_r_payload_data[511 : 480];
    end
  end

  assign _zz_when_MemoryEngine_l311_3 = (loadReqEntry_wordOff + 4'b0011);
  assign when_MemoryEngine_l311_48 = (_zz_when_MemoryEngine_l311_3 == 4'b0000);
  assign when_MemoryEngine_l311_49 = (_zz_when_MemoryEngine_l311_3 == 4'b0001);
  assign when_MemoryEngine_l311_50 = (_zz_when_MemoryEngine_l311_3 == 4'b0010);
  assign when_MemoryEngine_l311_51 = (_zz_when_MemoryEngine_l311_3 == 4'b0011);
  assign when_MemoryEngine_l311_52 = (_zz_when_MemoryEngine_l311_3 == 4'b0100);
  assign when_MemoryEngine_l311_53 = (_zz_when_MemoryEngine_l311_3 == 4'b0101);
  assign when_MemoryEngine_l311_54 = (_zz_when_MemoryEngine_l311_3 == 4'b0110);
  assign when_MemoryEngine_l311_55 = (_zz_when_MemoryEngine_l311_3 == 4'b0111);
  assign when_MemoryEngine_l311_56 = (_zz_when_MemoryEngine_l311_3 == 4'b1000);
  assign when_MemoryEngine_l311_57 = (_zz_when_MemoryEngine_l311_3 == 4'b1001);
  assign when_MemoryEngine_l311_58 = (_zz_when_MemoryEngine_l311_3 == 4'b1010);
  assign when_MemoryEngine_l311_59 = (_zz_when_MemoryEngine_l311_3 == 4'b1011);
  assign when_MemoryEngine_l311_60 = (_zz_when_MemoryEngine_l311_3 == 4'b1100);
  assign when_MemoryEngine_l311_61 = (_zz_when_MemoryEngine_l311_3 == 4'b1101);
  assign when_MemoryEngine_l311_62 = (_zz_when_MemoryEngine_l311_3 == 4'b1110);
  assign when_MemoryEngine_l311_63 = (_zz_when_MemoryEngine_l311_3 == 4'b1111);
  always @(*) begin
    _zz_io_vloadWriteReqs_0_4_payload_data = 32'h0;
    if(when_MemoryEngine_l311_64) begin
      _zz_io_vloadWriteReqs_0_4_payload_data = io_axiMaster_r_payload_data[31 : 0];
    end
    if(when_MemoryEngine_l311_65) begin
      _zz_io_vloadWriteReqs_0_4_payload_data = io_axiMaster_r_payload_data[63 : 32];
    end
    if(when_MemoryEngine_l311_66) begin
      _zz_io_vloadWriteReqs_0_4_payload_data = io_axiMaster_r_payload_data[95 : 64];
    end
    if(when_MemoryEngine_l311_67) begin
      _zz_io_vloadWriteReqs_0_4_payload_data = io_axiMaster_r_payload_data[127 : 96];
    end
    if(when_MemoryEngine_l311_68) begin
      _zz_io_vloadWriteReqs_0_4_payload_data = io_axiMaster_r_payload_data[159 : 128];
    end
    if(when_MemoryEngine_l311_69) begin
      _zz_io_vloadWriteReqs_0_4_payload_data = io_axiMaster_r_payload_data[191 : 160];
    end
    if(when_MemoryEngine_l311_70) begin
      _zz_io_vloadWriteReqs_0_4_payload_data = io_axiMaster_r_payload_data[223 : 192];
    end
    if(when_MemoryEngine_l311_71) begin
      _zz_io_vloadWriteReqs_0_4_payload_data = io_axiMaster_r_payload_data[255 : 224];
    end
    if(when_MemoryEngine_l311_72) begin
      _zz_io_vloadWriteReqs_0_4_payload_data = io_axiMaster_r_payload_data[287 : 256];
    end
    if(when_MemoryEngine_l311_73) begin
      _zz_io_vloadWriteReqs_0_4_payload_data = io_axiMaster_r_payload_data[319 : 288];
    end
    if(when_MemoryEngine_l311_74) begin
      _zz_io_vloadWriteReqs_0_4_payload_data = io_axiMaster_r_payload_data[351 : 320];
    end
    if(when_MemoryEngine_l311_75) begin
      _zz_io_vloadWriteReqs_0_4_payload_data = io_axiMaster_r_payload_data[383 : 352];
    end
    if(when_MemoryEngine_l311_76) begin
      _zz_io_vloadWriteReqs_0_4_payload_data = io_axiMaster_r_payload_data[415 : 384];
    end
    if(when_MemoryEngine_l311_77) begin
      _zz_io_vloadWriteReqs_0_4_payload_data = io_axiMaster_r_payload_data[447 : 416];
    end
    if(when_MemoryEngine_l311_78) begin
      _zz_io_vloadWriteReqs_0_4_payload_data = io_axiMaster_r_payload_data[479 : 448];
    end
    if(when_MemoryEngine_l311_79) begin
      _zz_io_vloadWriteReqs_0_4_payload_data = io_axiMaster_r_payload_data[511 : 480];
    end
  end

  assign _zz_when_MemoryEngine_l311_4 = (loadReqEntry_wordOff + 4'b0100);
  assign when_MemoryEngine_l311_64 = (_zz_when_MemoryEngine_l311_4 == 4'b0000);
  assign when_MemoryEngine_l311_65 = (_zz_when_MemoryEngine_l311_4 == 4'b0001);
  assign when_MemoryEngine_l311_66 = (_zz_when_MemoryEngine_l311_4 == 4'b0010);
  assign when_MemoryEngine_l311_67 = (_zz_when_MemoryEngine_l311_4 == 4'b0011);
  assign when_MemoryEngine_l311_68 = (_zz_when_MemoryEngine_l311_4 == 4'b0100);
  assign when_MemoryEngine_l311_69 = (_zz_when_MemoryEngine_l311_4 == 4'b0101);
  assign when_MemoryEngine_l311_70 = (_zz_when_MemoryEngine_l311_4 == 4'b0110);
  assign when_MemoryEngine_l311_71 = (_zz_when_MemoryEngine_l311_4 == 4'b0111);
  assign when_MemoryEngine_l311_72 = (_zz_when_MemoryEngine_l311_4 == 4'b1000);
  assign when_MemoryEngine_l311_73 = (_zz_when_MemoryEngine_l311_4 == 4'b1001);
  assign when_MemoryEngine_l311_74 = (_zz_when_MemoryEngine_l311_4 == 4'b1010);
  assign when_MemoryEngine_l311_75 = (_zz_when_MemoryEngine_l311_4 == 4'b1011);
  assign when_MemoryEngine_l311_76 = (_zz_when_MemoryEngine_l311_4 == 4'b1100);
  assign when_MemoryEngine_l311_77 = (_zz_when_MemoryEngine_l311_4 == 4'b1101);
  assign when_MemoryEngine_l311_78 = (_zz_when_MemoryEngine_l311_4 == 4'b1110);
  assign when_MemoryEngine_l311_79 = (_zz_when_MemoryEngine_l311_4 == 4'b1111);
  always @(*) begin
    _zz_io_vloadWriteReqs_0_5_payload_data = 32'h0;
    if(when_MemoryEngine_l311_80) begin
      _zz_io_vloadWriteReqs_0_5_payload_data = io_axiMaster_r_payload_data[31 : 0];
    end
    if(when_MemoryEngine_l311_81) begin
      _zz_io_vloadWriteReqs_0_5_payload_data = io_axiMaster_r_payload_data[63 : 32];
    end
    if(when_MemoryEngine_l311_82) begin
      _zz_io_vloadWriteReqs_0_5_payload_data = io_axiMaster_r_payload_data[95 : 64];
    end
    if(when_MemoryEngine_l311_83) begin
      _zz_io_vloadWriteReqs_0_5_payload_data = io_axiMaster_r_payload_data[127 : 96];
    end
    if(when_MemoryEngine_l311_84) begin
      _zz_io_vloadWriteReqs_0_5_payload_data = io_axiMaster_r_payload_data[159 : 128];
    end
    if(when_MemoryEngine_l311_85) begin
      _zz_io_vloadWriteReqs_0_5_payload_data = io_axiMaster_r_payload_data[191 : 160];
    end
    if(when_MemoryEngine_l311_86) begin
      _zz_io_vloadWriteReqs_0_5_payload_data = io_axiMaster_r_payload_data[223 : 192];
    end
    if(when_MemoryEngine_l311_87) begin
      _zz_io_vloadWriteReqs_0_5_payload_data = io_axiMaster_r_payload_data[255 : 224];
    end
    if(when_MemoryEngine_l311_88) begin
      _zz_io_vloadWriteReqs_0_5_payload_data = io_axiMaster_r_payload_data[287 : 256];
    end
    if(when_MemoryEngine_l311_89) begin
      _zz_io_vloadWriteReqs_0_5_payload_data = io_axiMaster_r_payload_data[319 : 288];
    end
    if(when_MemoryEngine_l311_90) begin
      _zz_io_vloadWriteReqs_0_5_payload_data = io_axiMaster_r_payload_data[351 : 320];
    end
    if(when_MemoryEngine_l311_91) begin
      _zz_io_vloadWriteReqs_0_5_payload_data = io_axiMaster_r_payload_data[383 : 352];
    end
    if(when_MemoryEngine_l311_92) begin
      _zz_io_vloadWriteReqs_0_5_payload_data = io_axiMaster_r_payload_data[415 : 384];
    end
    if(when_MemoryEngine_l311_93) begin
      _zz_io_vloadWriteReqs_0_5_payload_data = io_axiMaster_r_payload_data[447 : 416];
    end
    if(when_MemoryEngine_l311_94) begin
      _zz_io_vloadWriteReqs_0_5_payload_data = io_axiMaster_r_payload_data[479 : 448];
    end
    if(when_MemoryEngine_l311_95) begin
      _zz_io_vloadWriteReqs_0_5_payload_data = io_axiMaster_r_payload_data[511 : 480];
    end
  end

  assign _zz_when_MemoryEngine_l311_5 = (loadReqEntry_wordOff + 4'b0101);
  assign when_MemoryEngine_l311_80 = (_zz_when_MemoryEngine_l311_5 == 4'b0000);
  assign when_MemoryEngine_l311_81 = (_zz_when_MemoryEngine_l311_5 == 4'b0001);
  assign when_MemoryEngine_l311_82 = (_zz_when_MemoryEngine_l311_5 == 4'b0010);
  assign when_MemoryEngine_l311_83 = (_zz_when_MemoryEngine_l311_5 == 4'b0011);
  assign when_MemoryEngine_l311_84 = (_zz_when_MemoryEngine_l311_5 == 4'b0100);
  assign when_MemoryEngine_l311_85 = (_zz_when_MemoryEngine_l311_5 == 4'b0101);
  assign when_MemoryEngine_l311_86 = (_zz_when_MemoryEngine_l311_5 == 4'b0110);
  assign when_MemoryEngine_l311_87 = (_zz_when_MemoryEngine_l311_5 == 4'b0111);
  assign when_MemoryEngine_l311_88 = (_zz_when_MemoryEngine_l311_5 == 4'b1000);
  assign when_MemoryEngine_l311_89 = (_zz_when_MemoryEngine_l311_5 == 4'b1001);
  assign when_MemoryEngine_l311_90 = (_zz_when_MemoryEngine_l311_5 == 4'b1010);
  assign when_MemoryEngine_l311_91 = (_zz_when_MemoryEngine_l311_5 == 4'b1011);
  assign when_MemoryEngine_l311_92 = (_zz_when_MemoryEngine_l311_5 == 4'b1100);
  assign when_MemoryEngine_l311_93 = (_zz_when_MemoryEngine_l311_5 == 4'b1101);
  assign when_MemoryEngine_l311_94 = (_zz_when_MemoryEngine_l311_5 == 4'b1110);
  assign when_MemoryEngine_l311_95 = (_zz_when_MemoryEngine_l311_5 == 4'b1111);
  always @(*) begin
    _zz_io_vloadWriteReqs_0_6_payload_data = 32'h0;
    if(when_MemoryEngine_l311_96) begin
      _zz_io_vloadWriteReqs_0_6_payload_data = io_axiMaster_r_payload_data[31 : 0];
    end
    if(when_MemoryEngine_l311_97) begin
      _zz_io_vloadWriteReqs_0_6_payload_data = io_axiMaster_r_payload_data[63 : 32];
    end
    if(when_MemoryEngine_l311_98) begin
      _zz_io_vloadWriteReqs_0_6_payload_data = io_axiMaster_r_payload_data[95 : 64];
    end
    if(when_MemoryEngine_l311_99) begin
      _zz_io_vloadWriteReqs_0_6_payload_data = io_axiMaster_r_payload_data[127 : 96];
    end
    if(when_MemoryEngine_l311_100) begin
      _zz_io_vloadWriteReqs_0_6_payload_data = io_axiMaster_r_payload_data[159 : 128];
    end
    if(when_MemoryEngine_l311_101) begin
      _zz_io_vloadWriteReqs_0_6_payload_data = io_axiMaster_r_payload_data[191 : 160];
    end
    if(when_MemoryEngine_l311_102) begin
      _zz_io_vloadWriteReqs_0_6_payload_data = io_axiMaster_r_payload_data[223 : 192];
    end
    if(when_MemoryEngine_l311_103) begin
      _zz_io_vloadWriteReqs_0_6_payload_data = io_axiMaster_r_payload_data[255 : 224];
    end
    if(when_MemoryEngine_l311_104) begin
      _zz_io_vloadWriteReqs_0_6_payload_data = io_axiMaster_r_payload_data[287 : 256];
    end
    if(when_MemoryEngine_l311_105) begin
      _zz_io_vloadWriteReqs_0_6_payload_data = io_axiMaster_r_payload_data[319 : 288];
    end
    if(when_MemoryEngine_l311_106) begin
      _zz_io_vloadWriteReqs_0_6_payload_data = io_axiMaster_r_payload_data[351 : 320];
    end
    if(when_MemoryEngine_l311_107) begin
      _zz_io_vloadWriteReqs_0_6_payload_data = io_axiMaster_r_payload_data[383 : 352];
    end
    if(when_MemoryEngine_l311_108) begin
      _zz_io_vloadWriteReqs_0_6_payload_data = io_axiMaster_r_payload_data[415 : 384];
    end
    if(when_MemoryEngine_l311_109) begin
      _zz_io_vloadWriteReqs_0_6_payload_data = io_axiMaster_r_payload_data[447 : 416];
    end
    if(when_MemoryEngine_l311_110) begin
      _zz_io_vloadWriteReqs_0_6_payload_data = io_axiMaster_r_payload_data[479 : 448];
    end
    if(when_MemoryEngine_l311_111) begin
      _zz_io_vloadWriteReqs_0_6_payload_data = io_axiMaster_r_payload_data[511 : 480];
    end
  end

  assign _zz_when_MemoryEngine_l311_6 = (loadReqEntry_wordOff + 4'b0110);
  assign when_MemoryEngine_l311_96 = (_zz_when_MemoryEngine_l311_6 == 4'b0000);
  assign when_MemoryEngine_l311_97 = (_zz_when_MemoryEngine_l311_6 == 4'b0001);
  assign when_MemoryEngine_l311_98 = (_zz_when_MemoryEngine_l311_6 == 4'b0010);
  assign when_MemoryEngine_l311_99 = (_zz_when_MemoryEngine_l311_6 == 4'b0011);
  assign when_MemoryEngine_l311_100 = (_zz_when_MemoryEngine_l311_6 == 4'b0100);
  assign when_MemoryEngine_l311_101 = (_zz_when_MemoryEngine_l311_6 == 4'b0101);
  assign when_MemoryEngine_l311_102 = (_zz_when_MemoryEngine_l311_6 == 4'b0110);
  assign when_MemoryEngine_l311_103 = (_zz_when_MemoryEngine_l311_6 == 4'b0111);
  assign when_MemoryEngine_l311_104 = (_zz_when_MemoryEngine_l311_6 == 4'b1000);
  assign when_MemoryEngine_l311_105 = (_zz_when_MemoryEngine_l311_6 == 4'b1001);
  assign when_MemoryEngine_l311_106 = (_zz_when_MemoryEngine_l311_6 == 4'b1010);
  assign when_MemoryEngine_l311_107 = (_zz_when_MemoryEngine_l311_6 == 4'b1011);
  assign when_MemoryEngine_l311_108 = (_zz_when_MemoryEngine_l311_6 == 4'b1100);
  assign when_MemoryEngine_l311_109 = (_zz_when_MemoryEngine_l311_6 == 4'b1101);
  assign when_MemoryEngine_l311_110 = (_zz_when_MemoryEngine_l311_6 == 4'b1110);
  assign when_MemoryEngine_l311_111 = (_zz_when_MemoryEngine_l311_6 == 4'b1111);
  always @(*) begin
    _zz_io_vloadWriteReqs_0_7_payload_data = 32'h0;
    if(when_MemoryEngine_l311_112) begin
      _zz_io_vloadWriteReqs_0_7_payload_data = io_axiMaster_r_payload_data[31 : 0];
    end
    if(when_MemoryEngine_l311_113) begin
      _zz_io_vloadWriteReqs_0_7_payload_data = io_axiMaster_r_payload_data[63 : 32];
    end
    if(when_MemoryEngine_l311_114) begin
      _zz_io_vloadWriteReqs_0_7_payload_data = io_axiMaster_r_payload_data[95 : 64];
    end
    if(when_MemoryEngine_l311_115) begin
      _zz_io_vloadWriteReqs_0_7_payload_data = io_axiMaster_r_payload_data[127 : 96];
    end
    if(when_MemoryEngine_l311_116) begin
      _zz_io_vloadWriteReqs_0_7_payload_data = io_axiMaster_r_payload_data[159 : 128];
    end
    if(when_MemoryEngine_l311_117) begin
      _zz_io_vloadWriteReqs_0_7_payload_data = io_axiMaster_r_payload_data[191 : 160];
    end
    if(when_MemoryEngine_l311_118) begin
      _zz_io_vloadWriteReqs_0_7_payload_data = io_axiMaster_r_payload_data[223 : 192];
    end
    if(when_MemoryEngine_l311_119) begin
      _zz_io_vloadWriteReqs_0_7_payload_data = io_axiMaster_r_payload_data[255 : 224];
    end
    if(when_MemoryEngine_l311_120) begin
      _zz_io_vloadWriteReqs_0_7_payload_data = io_axiMaster_r_payload_data[287 : 256];
    end
    if(when_MemoryEngine_l311_121) begin
      _zz_io_vloadWriteReqs_0_7_payload_data = io_axiMaster_r_payload_data[319 : 288];
    end
    if(when_MemoryEngine_l311_122) begin
      _zz_io_vloadWriteReqs_0_7_payload_data = io_axiMaster_r_payload_data[351 : 320];
    end
    if(when_MemoryEngine_l311_123) begin
      _zz_io_vloadWriteReqs_0_7_payload_data = io_axiMaster_r_payload_data[383 : 352];
    end
    if(when_MemoryEngine_l311_124) begin
      _zz_io_vloadWriteReqs_0_7_payload_data = io_axiMaster_r_payload_data[415 : 384];
    end
    if(when_MemoryEngine_l311_125) begin
      _zz_io_vloadWriteReqs_0_7_payload_data = io_axiMaster_r_payload_data[447 : 416];
    end
    if(when_MemoryEngine_l311_126) begin
      _zz_io_vloadWriteReqs_0_7_payload_data = io_axiMaster_r_payload_data[479 : 448];
    end
    if(when_MemoryEngine_l311_127) begin
      _zz_io_vloadWriteReqs_0_7_payload_data = io_axiMaster_r_payload_data[511 : 480];
    end
  end

  assign _zz_when_MemoryEngine_l311_7 = (loadReqEntry_wordOff + 4'b0111);
  assign when_MemoryEngine_l311_112 = (_zz_when_MemoryEngine_l311_7 == 4'b0000);
  assign when_MemoryEngine_l311_113 = (_zz_when_MemoryEngine_l311_7 == 4'b0001);
  assign when_MemoryEngine_l311_114 = (_zz_when_MemoryEngine_l311_7 == 4'b0010);
  assign when_MemoryEngine_l311_115 = (_zz_when_MemoryEngine_l311_7 == 4'b0011);
  assign when_MemoryEngine_l311_116 = (_zz_when_MemoryEngine_l311_7 == 4'b0100);
  assign when_MemoryEngine_l311_117 = (_zz_when_MemoryEngine_l311_7 == 4'b0101);
  assign when_MemoryEngine_l311_118 = (_zz_when_MemoryEngine_l311_7 == 4'b0110);
  assign when_MemoryEngine_l311_119 = (_zz_when_MemoryEngine_l311_7 == 4'b0111);
  assign when_MemoryEngine_l311_120 = (_zz_when_MemoryEngine_l311_7 == 4'b1000);
  assign when_MemoryEngine_l311_121 = (_zz_when_MemoryEngine_l311_7 == 4'b1001);
  assign when_MemoryEngine_l311_122 = (_zz_when_MemoryEngine_l311_7 == 4'b1010);
  assign when_MemoryEngine_l311_123 = (_zz_when_MemoryEngine_l311_7 == 4'b1011);
  assign when_MemoryEngine_l311_124 = (_zz_when_MemoryEngine_l311_7 == 4'b1100);
  assign when_MemoryEngine_l311_125 = (_zz_when_MemoryEngine_l311_7 == 4'b1101);
  assign when_MemoryEngine_l311_126 = (_zz_when_MemoryEngine_l311_7 == 4'b1110);
  assign when_MemoryEngine_l311_127 = (_zz_when_MemoryEngine_l311_7 == 4'b1111);
  assign when_MemoryEngine_l340 = (! awAccepted);
  assign when_MemoryEngine_l341 = (! wAccepted);
  assign io_axiMaster_aw_fire = (io_axiMaster_aw_valid && io_axiMaster_aw_ready);
  assign io_axiMaster_w_fire = (io_axiMaster_w_valid && io_axiMaster_w_ready);
  assign when_MemoryEngine_l353 = ((io_axiMaster_aw_fire || awAccepted) && (io_axiMaster_w_fire || wAccepted));
  always @(posedge clk) begin
    if(reset) begin
      loadReqValid <= 1'b0;
      state <= MemState_IDLE;
      awAccepted <= 1'b0;
      wAccepted <= 1'b0;
    end else begin
      if(when_MemoryEngine_l180) begin
        loadReqValid <= 1'b1;
      end
      if(when_MemoryEngine_l285) begin
        loadReqValid <= 1'b0;
      end
      case(state)
        MemState_IDLE : begin
          if(storeReqFifo_io_pop_valid) begin
            awAccepted <= 1'b0;
            wAccepted <= 1'b0;
            state <= MemState_STORE_AW_W;
          end
        end
        MemState_STORE_AW_W : begin
          if(io_axiMaster_aw_fire) begin
            awAccepted <= 1'b1;
          end
          if(io_axiMaster_w_fire) begin
            wAccepted <= 1'b1;
          end
          if(when_MemoryEngine_l353) begin
            awAccepted <= 1'b0;
            wAccepted <= 1'b0;
            state <= MemState_STORE_B;
          end
        end
        default : begin
          if(io_axiMaster_b_valid) begin
            state <= MemState_IDLE;
          end
        end
      endcase
    end
  end

  always @(posedge clk) begin
    if(when_MemoryEngine_l180) begin
      loadReqEntry_slotIdx <= 1'b0;
      loadReqEntry_wordOff <= _zz_loadReqEntry_wordOff_1[3:0];
      loadReqEntry_isVector <= (io_loadSlots_0_opcode == 3'b011);
      case(io_loadSlots_0_opcode)
        3'b001 : begin
          loadReqEntry_axiAddr <= _zz_loadReqEntry_axiAddr_1;
          loadReqEntry_destAddr <= io_loadSlots_0_dest;
        end
        3'b010 : begin
          loadReqEntry_axiAddr <= (_zz_loadReqEntry_axiAddr_2 & (~ _zz_loadReqEntry_axiAddr));
          loadReqEntry_destAddr <= (io_loadSlots_0_dest + _zz_loadReqEntry_destAddr);
          loadReqEntry_wordOff <= _zz_loadReqEntry_wordOff_2[3:0];
        end
        3'b011 : begin
          loadReqEntry_axiAddr <= _zz_loadReqEntry_axiAddr_1;
          loadReqEntry_destAddr <= io_loadSlots_0_dest;
        end
        default : begin
        end
      endcase
    end
    case(state)
      MemState_IDLE : begin
        if(storeReqFifo_io_pop_valid) begin
          capStoreReq_axiAddr <= storeReqFifo_io_pop_payload_axiAddr;
          capStoreReq_wdata <= storeReqFifo_io_pop_payload_wdata;
          capStoreReq_wstrb <= storeReqFifo_io_pop_payload_wstrb;
        end
      end
      MemState_STORE_AW_W : begin
      end
      default : begin
      end
    endcase
  end


endmodule

module StreamFifo (
  input  wire          io_push_valid,
  output wire          io_push_ready,
  input  wire [31:0]   io_push_payload_axiAddr,
  input  wire [511:0]  io_push_payload_wdata,
  input  wire [63:0]   io_push_payload_wstrb,
  output wire          io_pop_valid,
  input  wire          io_pop_ready,
  output wire [31:0]   io_pop_payload_axiAddr,
  output wire [511:0]  io_pop_payload_wdata,
  output wire [63:0]   io_pop_payload_wstrb,
  input  wire          io_flush,
  output wire [3:0]    io_occupancy,
  output wire [3:0]    io_availability,
  input  wire          clk,
  input  wire          reset
);

  reg        [607:0]  logic_ram_spinal_port1;
  wire       [607:0]  _zz_logic_ram_port;
  reg                 _zz_1;
  wire                logic_ptr_doPush;
  wire                logic_ptr_doPop;
  wire                logic_ptr_full;
  wire                logic_ptr_empty;
  reg        [3:0]    logic_ptr_push;
  reg        [3:0]    logic_ptr_pop;
  wire       [3:0]    logic_ptr_occupancy;
  wire       [3:0]    logic_ptr_popOnIo;
  wire                when_Stream_l1248;
  reg                 logic_ptr_wentUp;
  wire                io_push_fire;
  wire                logic_push_onRam_write_valid;
  wire       [2:0]    logic_push_onRam_write_payload_address;
  wire       [31:0]   logic_push_onRam_write_payload_data_axiAddr;
  wire       [511:0]  logic_push_onRam_write_payload_data_wdata;
  wire       [63:0]   logic_push_onRam_write_payload_data_wstrb;
  wire                logic_pop_addressGen_valid;
  reg                 logic_pop_addressGen_ready;
  wire       [2:0]    logic_pop_addressGen_payload;
  wire                logic_pop_addressGen_fire;
  wire                logic_pop_sync_readArbitation_valid;
  wire                logic_pop_sync_readArbitation_ready;
  wire       [2:0]    logic_pop_sync_readArbitation_payload;
  reg                 logic_pop_addressGen_rValid;
  reg        [2:0]    logic_pop_addressGen_rData;
  wire                when_Stream_l375;
  wire                logic_pop_sync_readPort_cmd_valid;
  wire       [2:0]    logic_pop_sync_readPort_cmd_payload;
  wire       [31:0]   logic_pop_sync_readPort_rsp_axiAddr;
  wire       [511:0]  logic_pop_sync_readPort_rsp_wdata;
  wire       [63:0]   logic_pop_sync_readPort_rsp_wstrb;
  wire       [607:0]  _zz_logic_pop_sync_readPort_rsp_axiAddr;
  wire                logic_pop_sync_readArbitation_translated_valid;
  wire                logic_pop_sync_readArbitation_translated_ready;
  wire       [31:0]   logic_pop_sync_readArbitation_translated_payload_axiAddr;
  wire       [511:0]  logic_pop_sync_readArbitation_translated_payload_wdata;
  wire       [63:0]   logic_pop_sync_readArbitation_translated_payload_wstrb;
  wire                logic_pop_sync_readArbitation_fire;
  reg        [3:0]    logic_pop_sync_popReg;
  reg [607:0] logic_ram [0:7];

  assign _zz_logic_ram_port = {logic_push_onRam_write_payload_data_wstrb,{logic_push_onRam_write_payload_data_wdata,logic_push_onRam_write_payload_data_axiAddr}};
  always @(posedge clk) begin
    if(_zz_1) begin
      logic_ram[logic_push_onRam_write_payload_address] <= _zz_logic_ram_port;
    end
  end

  always @(posedge clk) begin
    if(logic_pop_sync_readPort_cmd_valid) begin
      logic_ram_spinal_port1 <= logic_ram[logic_pop_sync_readPort_cmd_payload];
    end
  end

  always @(*) begin
    _zz_1 = 1'b0;
    if(logic_push_onRam_write_valid) begin
      _zz_1 = 1'b1;
    end
  end

  assign when_Stream_l1248 = (logic_ptr_doPush != logic_ptr_doPop);
  assign logic_ptr_full = (((logic_ptr_push ^ logic_ptr_popOnIo) ^ 4'b1000) == 4'b0000);
  assign logic_ptr_empty = (logic_ptr_push == logic_ptr_pop);
  assign logic_ptr_occupancy = (logic_ptr_push - logic_ptr_popOnIo);
  assign io_push_ready = (! logic_ptr_full);
  assign io_push_fire = (io_push_valid && io_push_ready);
  assign logic_ptr_doPush = io_push_fire;
  assign logic_push_onRam_write_valid = io_push_fire;
  assign logic_push_onRam_write_payload_address = logic_ptr_push[2:0];
  assign logic_push_onRam_write_payload_data_axiAddr = io_push_payload_axiAddr;
  assign logic_push_onRam_write_payload_data_wdata = io_push_payload_wdata;
  assign logic_push_onRam_write_payload_data_wstrb = io_push_payload_wstrb;
  assign logic_pop_addressGen_valid = (! logic_ptr_empty);
  assign logic_pop_addressGen_payload = logic_ptr_pop[2:0];
  assign logic_pop_addressGen_fire = (logic_pop_addressGen_valid && logic_pop_addressGen_ready);
  assign logic_ptr_doPop = logic_pop_addressGen_fire;
  always @(*) begin
    logic_pop_addressGen_ready = logic_pop_sync_readArbitation_ready;
    if(when_Stream_l375) begin
      logic_pop_addressGen_ready = 1'b1;
    end
  end

  assign when_Stream_l375 = (! logic_pop_sync_readArbitation_valid);
  assign logic_pop_sync_readArbitation_valid = logic_pop_addressGen_rValid;
  assign logic_pop_sync_readArbitation_payload = logic_pop_addressGen_rData;
  assign _zz_logic_pop_sync_readPort_rsp_axiAddr = logic_ram_spinal_port1;
  assign logic_pop_sync_readPort_rsp_axiAddr = _zz_logic_pop_sync_readPort_rsp_axiAddr[31 : 0];
  assign logic_pop_sync_readPort_rsp_wdata = _zz_logic_pop_sync_readPort_rsp_axiAddr[543 : 32];
  assign logic_pop_sync_readPort_rsp_wstrb = _zz_logic_pop_sync_readPort_rsp_axiAddr[607 : 544];
  assign logic_pop_sync_readPort_cmd_valid = logic_pop_addressGen_fire;
  assign logic_pop_sync_readPort_cmd_payload = logic_pop_addressGen_payload;
  assign logic_pop_sync_readArbitation_translated_valid = logic_pop_sync_readArbitation_valid;
  assign logic_pop_sync_readArbitation_ready = logic_pop_sync_readArbitation_translated_ready;
  assign logic_pop_sync_readArbitation_translated_payload_axiAddr = logic_pop_sync_readPort_rsp_axiAddr;
  assign logic_pop_sync_readArbitation_translated_payload_wdata = logic_pop_sync_readPort_rsp_wdata;
  assign logic_pop_sync_readArbitation_translated_payload_wstrb = logic_pop_sync_readPort_rsp_wstrb;
  assign io_pop_valid = logic_pop_sync_readArbitation_translated_valid;
  assign logic_pop_sync_readArbitation_translated_ready = io_pop_ready;
  assign io_pop_payload_axiAddr = logic_pop_sync_readArbitation_translated_payload_axiAddr;
  assign io_pop_payload_wdata = logic_pop_sync_readArbitation_translated_payload_wdata;
  assign io_pop_payload_wstrb = logic_pop_sync_readArbitation_translated_payload_wstrb;
  assign logic_pop_sync_readArbitation_fire = (logic_pop_sync_readArbitation_valid && logic_pop_sync_readArbitation_ready);
  assign logic_ptr_popOnIo = logic_pop_sync_popReg;
  assign io_occupancy = logic_ptr_occupancy;
  assign io_availability = (4'b1000 - logic_ptr_occupancy);
  always @(posedge clk) begin
    if(reset) begin
      logic_ptr_push <= 4'b0000;
      logic_ptr_pop <= 4'b0000;
      logic_ptr_wentUp <= 1'b0;
      logic_pop_addressGen_rValid <= 1'b0;
      logic_pop_sync_popReg <= 4'b0000;
    end else begin
      if(when_Stream_l1248) begin
        logic_ptr_wentUp <= logic_ptr_doPush;
      end
      if(io_flush) begin
        logic_ptr_wentUp <= 1'b0;
      end
      if(logic_ptr_doPush) begin
        logic_ptr_push <= (logic_ptr_push + 4'b0001);
      end
      if(logic_ptr_doPop) begin
        logic_ptr_pop <= (logic_ptr_pop + 4'b0001);
      end
      if(io_flush) begin
        logic_ptr_push <= 4'b0000;
        logic_ptr_pop <= 4'b0000;
      end
      if(logic_pop_addressGen_ready) begin
        logic_pop_addressGen_rValid <= logic_pop_addressGen_valid;
      end
      if(io_flush) begin
        logic_pop_addressGen_rValid <= 1'b0;
      end
      if(logic_pop_sync_readArbitation_fire) begin
        logic_pop_sync_popReg <= logic_ptr_pop;
      end
      if(io_flush) begin
        logic_pop_sync_popReg <= 4'b0000;
      end
    end
  end

  always @(posedge clk) begin
    if(logic_pop_addressGen_ready) begin
      logic_pop_addressGen_rData <= logic_pop_addressGen_payload;
    end
  end


endmodule
